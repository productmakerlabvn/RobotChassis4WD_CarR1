PK   �A�X�2#�  ��     cirkitFile.json�][��6��+��.`yx��[.l�I#�]�%Q)o�v�lw'�����|�-�>�a�l:A�,��G��s��yT��~�X,j������b>��r<zru�ɵ���y:\-������s���~�Y������Q2�8*��2�D�ifh~JE���B��������)�9�5��"4�k̉�N�4Ӻ��`LgF;��x��e�#z�8��q�a\�7��	V,ؑh�H�S$ީ@�G*d{$�(~�?���J[$�lH�:�{�s�UJ�L�f��y�9�5S�iZD�a������!y뛣�֨�Qʂ�����t�q�\�|x���<�/K���e��e&*Ufy�eF|���E�
��ގ/-a��"��gF�:c�)��sɼ#���	��!;�5�Zx�LY�FdB�И���s�d>7����☞Q�<lD���ak�tA2N�΄aE�H(��I�9�n�ZsQZ�3R���S>s��S.�\0�[��!	�z � �QS���������yH�äj��腵V���(p�0]IA����{HB3L�C�,� ��=$F��8�o�9;$��:�5�Å&�:��F3�Cfs"2�+啢�SfP{ �-�k��zH����a; C t����!� t0�rH
�%L�C���pX��^��.�0��&!B"AhB#z�Y@������x�5�3�3}��Q�<4�@G�t�p���~_�X�5r_m�7�������TX*<	�T��LJBE'�b�P�iP��i�K�����/iȤA0Ma��4�i�4(f�dp�4(f[ˊ[���^���?��p^�V��o�b<�L�ₙ�V2[;�1��4(�Q�[
#���A�nP���m@�^�[�}��rQ)@�FFS��<GPQ�qa�DP٬%Z�ËIB�YIȄ;��f`,Z��@{
n�%a����P�yA�J�W+� ����Ɗ�h���҆�RP���M���ޠQ���<�D�8��х�������X�y��۝W���y���%�B/=4�u~t�1��L�O˕[yl�i�׫�͐�'<��
OBE$�"�PQI��$TL*6��7zi��4��i L� ���0M�a��4�Y�D28�Y�4(fiP�Ҡ��A1K�b��<��E��Ox*ix�����'<���	�S�����'<��K	J��D�M���V<���L _�j��d��'<����?ᩤ��"���'<���ǟ�Rǟ�T.�8���r�p�	O�"/����E^��'<�6/_����&��qZ�6��v<�4����y�
_>N珋������J���4�L|T�AK�a�V����[�|EL߯	5�f0�M�FY͘�1���5���y���h���1������~3�\
�x6*,��%D��l��4`z�$eᄷB����4���s�|b �����y�{���(��>˞|UAϣ��y����\7/���w��׳����Q'�1��{�jоJ�.K��K���$�7Xw�ҫA�l�)Dһ�3�t�� }���.���u��?��s���� �1<H�������v��?�U�3����S�t�%8���@u�^l����Ϲ�\O������E�Mˏ9��i��H~D�"c�3d{�l�����{'��.;����d{�E�X|R,@)�M� �M�� �D�E"�"��%%��D���t�.=��z��'�P��MW����.�p,����3�Oh�����0���'Í	>�.9L錚 ��ր?N8>!�y�@�R� ��Q�z"f�hwpiw!���Y	(��g)�Ο�C��?��3�QT��i>!7 ����'�8�y@0��O�10��D�rXg<�ր�>�p�y����C8�,p>��`,Kpb�	�)	ΐ>!7�c���'�d8g:!��0!����N�ʗ��@fZ�`Z����4���j�fQE�E�(�G��$�;J�f7b�]J�jƼ)��؀�,�`�؂�,�`��-Xl�b[�؂7o'�(���>!�������e�5�d  �8G=B��QȺ<j Y*G �m5�]o�:�����K�Od*����T��)���2;�k	�9�L�����o!s��~�ȴ��U���2ӿ�#�>݂K��b�7�c� ����	�z�;&�K����ϛ!��~�;oȔ�����:*.˾�?��1�K��Z��b�G�QwdHu`>"��$mw!��0N.�낡>7�qQ(;wO����h����%�ӯ�"�'%t[D�El[ĺE|[ĻEb[$�Er[$�Ej[��Ez[��Ef[d�Ev[d;Et7�;t?������������!��!��1��1	a��l���ޕ����B�x�M���\��/�p����Te��2�	�������G����-�`�<f�<���b ����/�u���}nn��Ͼ^M}��<��D���z:�%<��}��c�x������W�d�Y^ϧ��Q�Z>->�0�&��W��P������4������k=�}9�_�kF䃛�+W�ֵ��1Ю��d�$�������r�j>n�NI:ar��D��L�	5G����gZJ�iA�pgyfr�h����ڏ�Ͼ^6�x4�/Wn^l�b.�Ѣ�*n��(Lt�=������;��ca��Їkպ�[���&�������}պ6�:�p���}�Z����&\3B���kE�k����u_���}{������Y�ג�U�iݷ�����^��}���,�2QJ6������hF���~U<=���i�ܑԊ<7UV��D��g�W2ӄ˲�T(�������"���Vfo6m��J� ���/nx�(�2bi��p�(U�6��jg�־p6�}^�>�"�U@��I�h*�վݛ��z�j\��_��"������V�<׎�\����#��Ø<���I�y���� �HP�6�eP�B�<sU(sf���Ɉ������b�ó������0�EX�J���e��"�i���ˈ+{�|3[,}�Uh^X����	���*(~W�������s��g7/}leG��MV�:������7ӵ�y�>�����iܮ��J�%o�ꫲ��r�-�2�c�Q5��pM�[�[�y�-���?2�a�Kg�h]p��C 3��B����`CV<SƗ�	z�p�`�o��R��2����3�̌p��d�-fu�R�D\ܰ"B�+�J���ک�T�Vl~>�>.���ү����w��ww��]����źޔ���wO�����^��A*߇���/�B�Ţ��7������w+_�~o�p����b�@���˘�G�����{��=4��(���~Z���b�LFt�'1��U�����l6�_[��ݏ�|�J�ȕ�Ha�5r�I9RI#��k�v]Te&�s�P�VY��לs_Y�j�G T�l�L���\�IPL���o�)�h���c��F�32ђkJO��"Bؓmi��
KC��������'�0����h��&���d"b����l���n�0����C&�0�j��`>P����-.c1e���֜I9vC(�l�Mc(4���Śn:g���mZ�]���DC�
�_|x�n�y�̟`�U��^OWwo��:�	�z�0�F��e��Uc!Ʉ2}���w�;n�^�,(���QO�a�
_�e!��������z��Ӫ���Ʋo������E�N���H���1�Ԉ	��4��uʹ��u2��.�dE(��F�dF��:���.��!��eD��l������C�KT�D�� ��8y�5�����kR�1WGk/.����a�x[��?���9��jI@@���W����5�mi]���:���)����]��w�y�駄�	T�D�gTN�`J�	چ����12�x48{YY�2+�Yn-�0����m"+'�F�a��>h��e	c{��/ � P��$X�B�L�`Frj�ä9���F��@�1� *���&��F��&�H��Ẹi��fg����4��[�Y�
��(;
����<�8,j'}8��XN��;�V���D*�oE��M�a�%�}���@���8�Ǜ�m	�N$�EŽ��z^6�Y-�P��?��G��|�#�1�;ŗw���H"�H!��^ѓo�p��C��N��~�ALluœ/��o����j���S���K�����%�-�&L���a��]��N��`�����<K���Ъݧ��2�#!ϋ�|�֭�b�Fq���m,��Y��x��]���e�6c�qO-z$���A�+j�c-r[����ї �cll>d�*!6xjl����7a#��]��q��Y?D�����I�!bC�ƆL�q6$HnH��8�o%�Tn4��M��256DZlț��Ar����>hE- 66�jb�?��kxK{2Z�@��4�ԋ��vW�oL]R'���IaA��$��P�����[�L�{*AWy���әЩ0�'3�KanZ����f��v�+�R�L8T:�J�+�w�ϭ���,�@q��yk�@q���������~.ّ֢��V+^�w�D�t�k��
��D��Ŏ��N�!o#50�W�(�`-�X�)Bq
��܋�drrS�^uÌ������C*�PD�a�_�Wp�"H�Rk��=Q�ZC�p������<C
G���q{WBc��t�� ���vK��a�����~��J�!XLx�71��!�k��bH��'%'�7X�#�9usm-(���	1��a������M���4��c`5Ib�G}�j	�dWya�S��tŦ���B�M[>�u$t��$���c�j]�������
!��v����T��M2Ȫ���5I��_H��C/-Ŵ;3P+(`�xP\�ګ���贙�}��<;��j)��/9t/�ʑtظb/�
�Ra㦝�V�v�J`���z�
���ё�A|�VJ /؛e^^W�����$`��E�.��~2���� T)%ʪJǓ�o�P{�P��m(ʮ��J�ɣ~��G3)�����E�`��� �>=0�x�`o�J'Į�<�YK�;q�Z'U�i:V9R����:P�^ ^ �@�2Λ�R��`�
K,u���
�pRg`�sC�~���c�R��xLK�Y}�J	 {	\:�sͦ<��Tr�&���k����)���x�hĳ/����{����͖����e�c�o_~��k7�z�������y�>"�^��/V��eQO��gwF_�PK   �A�X��_�  >  /   images/17d126d1-8a97-48c5-9cdb-beb53ba7b71c.png�XgPP���:�PZ�� �*"U@@z $*B���ބЃH/�� �{���ޔ�q3��~�����̾�y�;�����}1&F��@
<<<j]M�;�|�cd$w�Qs��!�ձB��qu������?��dCjY"�<G8������<N��.b>~�Y�J���!]Mu���=���v�/�����z[��l��։�Ll��BHJKu�9P��	�P~ۻw�����&2��D Xj���=í��¼�E��D���(���\��l�_4�(U�qOؿQ���;r�s������@u�$
��P��a׈~�KfJE��i���3���tL�OO~�����~��.L���(�,x�����Gy-�Ō�*��4�RϿ''�����42b�j�����-�<��v��ZJF��>4z��/��z�F�8\7d�&���>���ؼ�����		/���s���@<�fa#��	����09�z���ڵ�P��lI����a��>sO���72=1��SI�Y��'���哜i
~(�#Z�pG�<\���ssr��`�����B�)��(΅�����Hj��Rrޓx"S ��Y��]:��CΗE5�V���m-�"�ǵp���eD_Oh���\��V��B�����I"��u�X�i藻e#��D\�(�d�s�I1��]^Η�N��v�0�h8 )�37�+q�o�F�U��x��Z<��W0�\; d�ھ:�m�gN.�+��R=r�c����MZ �	��3Go1j�֩��}0Ä�"��h<\�IO�뱀�"[/��'G_�Oj�t��������u����J�s9�੣�2���]D{^������i|L�M��eW%��w�2�
���0O����߷�qZ[�B��,��@�Ǭ��ۺ�{mG�k,��0ZA����S~e���X��p��d��
]]y M��1^?Ν���e�e����:t�w��ۋ�5�ψJ7�N��՟юmB�A&%�$�4Z���Qe|$2 n���9�Wmw�����[��S���%�z~�9�T����#����W������ɽ{X3�p��1�j�I5}J�'�*���X�9��FFZ��ɓ��J�0ż|�̎��G� �^���j��O5^�z��iz^���Ky'k��bYJUю?�f9ϑu�����2$�busK��=(�|��n+��*�u�R���񎔀��w�_s�b��#d�?	\l.+��1IO5�ɶ�`OP�(��^��eM%,?�������=�i��b�(��P<kk����ż���`�	o/�Umqnŋ�_\�iq췪���b�yh���\���][;)�9S^T��k�J���$��jo�r#if�fNj��.��N*<� 7KK1�N��V�d���,�CZ�,�es�iDԷ���EV�~��C�s��3,�,x�Q4[a�mg�W���@IA
���Gޢ<��w����i'\}}�0_ϭ��?�p聈�R `�Ǐ���F�PPo~\�2�B����d�.�	�
|-���I�H˖C�)�wl�9��zwӼ��_Yy����c�ZsV�dn��530�dtv��8��"�:ZZ2�0��r34ig*p��&����e���3�Z�"0k5.�+���IР<-Н67]"��Ȗ����z�8m��eD���[� ZJ��F��y�>+=\3')�_�(�H�9:	�iɉ�18����"2����=
�t��G|�(lc�Ÿ���A�����s<��<����e��z��Ht>�MJ�!�-�CL$߱���G�;��vӰ}B�'���#�"jY_1��X$�ˈ��ω�U��Y֔�I#s�nAl�($J���ޣ��i!�#	Jm���h���j<�Kg�Tɮ^������������*0g�������'���_O��
�6�ҥ��i�>����5 �\վӏ��Kz��ZH4x�h~�s<!i�F$.��#w��;nO��h��4xG����^�o��a�����\�/��EDN�q����$��~QqE���4�&����⧳�RQ$�ҹ����\o�r)�P���4[.���HR���Ie�h�g����J����g1M�В�hK^Á�kG�7�����)s�������-=O�<Ɖ�^d\��.N���u�0�iݲ����`ε?�8��*1/�o�?A'�p��a���	�vV@���\}�$o��������K��\���B���`��ɐ2����ᗰ,�*�ow�u�uT�c�RA �M�e$�2yt�l4��Q�͏�~�>���R9���kU�^*��xλ(�;��z����vf)"㕫�g<�������ϟ������i�G��#�F.�%t;"����v��k5�EE$%$$�$�@��nS��f���e�M���ө�ѹ���gTvڒQ���=r�&Gt^�3��s(��ok��͆�R�Z��,�1���,���B�KYo����2����|L�l���U�[^��O^����
�����2`�Dy�0rQ*%��y�Fs�K�`v9��/��MLL����P��3������͛���)�v�P��)����>XCDȇ�P���i��'?:��z��Yu�����Vz;~\�D��1|��o�s�4�z����3'�D�Ga�/څ�g��~P)[v){��!ejjj_�GWf��ﲯsY���%�'��_hSnN��7�+���$�ak�
?����<l{#WG=<<b�Z���;�IgcY+�O�W������o|T������o\U�JG���pW�~{�Dbv-���F�	U-zf{�|a�/����+�3W�<Tm�p5Bm���-�[�F�Tra=8�/�%���}�nT��^4g�i�L�8���h7Br��)���B��ާ�ϷV�5 H�}��B���q�
���-Թhj��7Kv������
�S�^��	�!r�<Y�\ �֑ �\�x
++��Ly��ց:]-�8}��F�i�`Q�ilg��˲b�{k����>��C��>����%����2��k%�:�賋����V<mm��g�ƒ���J��h͒,��h��"4�� �P]�(������>�}�'>?���ٙ�J��	�o4˳���{�v� �rl8�A�$����-�,�]����(��T{�_�����NOK��ėj��p����3���]�d����fP'8���Mn����&��"#EoD`D��B�Q<"3���$[D��a��^�S��eïI�ES��y�����\x�Ѕ#����^�
���O�,Я��@&_ ���9z�G�-He��恔'���]Mm���JϪq��^�2�yJ8f��SI�+��XHN�PD�-=���o��v�"ڋL��I�A�c��JKu���0(~*��,[�G����
v�:�?�p*�T`��dwpz��o#���IM#D� �C��y��,G�A�b�QR��D�M�2��&J�����C�� �:�>jn����=T�DD���&kYiW��	d��AXe���k��`>o+ATO�_OTĳ�|�`��(�S�)6��$�1�T/aً�,��$��K�浨��X�e�L�j�é��x�[+���V�@��1���p=����&�S�B�z|�N��ږ�J�YL�?���J���!�A?)EV��+HLo\��'2�f]e�4(ZL�;��0�|�q$R0_���GN�9#Z���"?QGf�7ǉ�+�O�+D�o|�/Ҋ�W�N�p�2`�X��~ֹ�&�y3�U\��Ա+�w��D�6�-�!H���k�>��/��V���АK�۝-���j�J�>�Ւl����s��������ݷk}b�v]W<��}�يo�K��&�W֑�1 ��<����/��Q܆�=|�ID�a#<<��7ZL�1 üTFg�*��75�f��p7����5븥��a���˵����q�ڢkT�y�ۇ��M�-A�c���g�D1Ѥu?6=��ϱ���\��L<����ֲw��
,��l�G0�M�j��/��ޙO04��('}��F���h��j2�Fpǘ:X�L��'�]V��NN�%�&����	k0�&��u��}��wA�}��\{�����f�do�F��A�j�RbC�&5b3I���R	c���himݙ�hݩ/�A�,��S�X	F|`@��nH�3��_�L��2/۸��%����v[-�?�Zݟ�&zapj��$͘m�!{�M���l�������{�?�$;I�x�oh�.
u�7�!���Ѥ�b'|s�zg�-�e�H:`A�^����bk�u<�꟢1�,�볤�s�0�P���W����^��Pi91����_�g��m�X͎|8�}��L/x�(Ј�����A{w�~��5�N��Yv"w;���>e�(��Ũ|6�h��(`	��W��s��|z"Q&$��|I�CqR#���W��C�cYcھpw־�ϛ����O&o�٫���k�k����7ׂ�c������F�}_�<J|6n�ls�C|�hW���e�]�	TT���$-�!�3+�r�ez�8��8�3��ۙ����7��c����'�ܞ��� BP��;2d`�	����<�Y��8U��vt�n!���#I.���I�u��H(ueY{��k#�X��|�5�9|��y����P��>
G�U1"�E6��Y7�~�IP�� lBy6'�T�m��Ҹ�}&^�BD
��#�d�_p4	��{��� �>۔�o��렡��������+C7��س�?�q�/�O<K&ʷ�	�)����*;�.�q�aD�ב���~�K����q�o�rF�Nܣ�Vsx��XH��������?�����`�s��%]�~t�U�y#�磪Q�Fn��!A����!�x��=�)ɛ��dee���2�9�+ �����W��'�fzqV�.��j_:�6�Cɜ�&�[n3ע<�S�P��d;�0+v�M֥��9��>?�8Ra�TЎc\�����M�3��vH(	�������dy�>��R�u#��&Ʊ���F�8���%�t����l�^6;�4C�@�-�^A�4�����?`0�XY��ʡ~����@~Cߔ7[b:��գϻY4�{����+��{w�Xgz��D� �x��K��������^��h\�[QCC�a����0���sħ,ߌ:��h!>�^��:6��"��*�,1�<��P9�.951Q�iiiѥ��i�X�ǙW�y�I��>-��g��nJ=��Z�����t����AX��W<�kA��*����l=���� �	4�ި!�$^�3'E>zN���MP{Eu{&�����ґ�_l�ߓ�����,���b���E��|����$i? qU��H�[�#��z���'�'��U� ��n�T��rx��l�O2EmV�SQk�$)�����A�~7����Q[i{�U�0��&��5ʖ+`�S�遇���ۨ�6��ɎZ����Uq�
W۪��N�PN3��'�8��I��������)�>[�x��*ب��i�}�V�vK�5�qM��{cr��Ud ��)�^끕^�'��i'b�ӥ�� ]J�F$�tn���o�t���b'�.��Ï��%1���c"�O�K:�J�/�<��o �� ��\-^2�7��)���%�Ա.K��ՓW������*j;����m=�N�jGI$ɇ�tY��uf�J:�(V���*��'�b&�̈́�s�NN$e��9[e��J��R,=2e7��lË�T��T}��N��U��>i5�1+��W�X��Zu˿�\���ն��"�c?
Oq���^�|n�~qz�؁�ӛUUu�0/�Ԭ�``=G�#_u��E�֝AZk���8�&�O�6L�a5��'��%R#����s�;�8Vx�-�%��V�J������V8��i'���ȹ!�*S}�`�1�WM<|r�9~����rTYq��A�,q8��j1�G@p���W�;��o /�4C^�����8;p�!���W���C�Oo�REӵ�}ձx[�o�LI��;U��ə7ޜ�.�f?�C����Ozi4>����>�.�XhL��|���V�n�nWf�l6���Ǐ��ӈ�#���z(�ǚtݝ��E�E
IYeq.DYC*��F50婻b:22t��ITi[K�t�ƹ�}�tFdYt��j�"<j�g��#���5U��}6����ӂGR��τ�����ʭNx'�,��.���$F�tV4���Ә2h17�D�Q��ΑY������t~���������-�A�{�x���u���T��q7��S��ˢ���t�����W
0Ƃlf�G:���/Z*x�:�!��_^��\�u�I�)��{���� <�;�"�lɺd3��$�"��>zf0<:�+�]���<ARwPDR��&�$�l�����OHiD�o<���xw��e���8��PK   �A�X�K��]r  ��  /   images/2ad7430d-0d07-4e15-a76a-a5ad941878d2.png�wT���?�>(ՁQD)b�p��JU����|�H� *Ma��	iB�� � !�H��{�8󾿵�k�?�Z��w����y���>{�ޟ}x�<���p��b?�`�}\�3�����`�rw� #?�+�߶\���.���.����ʭ L�������u0x4P�f�u���;�ΰ��%wo� �;��J>��)Kp1����o��.��=�@n���Yށ�Fvߺ����qӗ��0;<�W�Rfb��s��'J��]0Z������I����o���$�L�˚^,�-7�Hj���;�;�ʳm%�w��U���3űj�7ޮ/U�5��#�+#�`�~Y^��A�ٛ!���q��y=G�d�M�Xoj3T[
�
��i8����d'�,1-�XXpk���Z,����p�}+OGrW���j?�����ܷ��>Yr��2<KChcU��Z쾚i��!{O���w���6H
~���<�������@���ׯ_O�ϫ)�; l#�Ҭ+�ݖ�X��0��Y7J���(�y@�ag�?���]��5���4\�O$�O���Q���[/��Q�\����$���k�'��索�������瓹	���������m!7mz�%��}�3�$)�~�ڨp7��7�핝b��k{������!�MD�IM3�nе�q����H�y�|6k:Շ�L�	|u��P�I4E��9�����#q��Z�N�,.V������t=ʭ�
�����yy2�}�:�#	G��iL�79���i�Fkq�!/^��Ǐqb��E?x�`��� dS˄���j�k�{{��6�G��_�Sٺu����=z}�r��%� �O�^��+p�/� �~Y��n�O��Z����)4T�ɓ'E�mk����n��ǻ��3�z��_OՅ@k��hS�9��YK��6��9#�U�J�������������w�nM==��ʊe��X�B(d�������s��
�������Z�P��Д�i�;w:yy) Ų�i+|ՔΛ����7o�DgggY�+ ���j
dt�	a��#��K�~��'8��-����"�eC�̗))�ۃ��ܵ��'m�Hog����%�O$����SSS*gϮ��0�	���,�(�f��6H�g���JkFr֕��;��ه���TTT��R5���iiq�^�Jތ������rg-���p���b���'��e<ʇ�Y]*ZZ�d|fccÂ�,H"5�B���H��/_����%š�u��QL:����Kt^�R�C�����R�|H�[$�> �z�TQ�2�,Rn^��a�5=��ϗR��Uggg-�/F�^�����;Ur**{�+rٟ$.-��W�?4�:w� ��`p���Ќo����i�D��8�Ğkʬ�������u����N����X�H޽�|�^=�+�߄�ӫ��5V�\�\#��էr}�(㗯_���D��0�FBT�IQ�W3�����Y=hᆂ�B��� /��T]N~�kf��=7�Q(1�6�-߾}�>g ە�q���WrHN��Ͷ�І��FcfR�7� 3���&�k�9A� ���~}妚"9�(��-���
� �H1�J���B�M_�<�*+*6�Ecbb�O�4n)
�
^�na��	�e��ʖ8w�����h}u�ur�:��o�(("i��]iZ�߲W��U�s��jޱ�����
�:nd�a+���m��Z��Tz���i��Ɂ�I/`�Je�$���ե��d'�6nXX�i�g��RW��ʧy����%�녠�)���h��{Ӷ"�w]p��X�6hjU
���=Sq�(�D*s)�n�'��T��%�*�[��g�w	YY��vmܶ�����N95X �6wc|����7m��xW��k׮q=�"��բ������,,<���Tґ�!�;����[����F�)B�?'J
�~�zm� W|����r��Ԝ�Zkk����Ys��g�a+w�%e U���69��F�ה#�1�����w-�\�&��O�b��][�kpa�Y�oq���T��G�s�Dte��-���u"֛K��tp�Z䆩�Z���Qr,զ���>qՏE)�.��~2 �4+���dx��8��e뇩������ƲL0h!�@���� ������88�빒���6�
�g�I ϐ�V���y���}߻}�X��ce�e���� Ng�.�睊 w�$�u	:��єb�Γ�(�5�vz��w��Ff��0^b#���|7����wD\��TE�tgN����5�y���*1�* X���J�d=����?5�sKM*���'��Z�%G�L5�����AyD�G�B��AZ���E�!�ه��k�U(+)����{�#�6hRڈUJ���>'M}]G��ȣ���>,�_�\� ���5=lV�D0���B��<A�f
HO����$�����;z{+H�R���W�@�p�@V$� Uɜn�XG-hJ�n:Xkκ[6�A�L�0�Av�x�����<ߘ����:a����$��Ue�7@,��('~�s�6d�x_�}q+}�U�0��9���=#`:��UeJ���2�#FHH�u�3�f �2��d�H��D#i��Q�Cv/��mp��2����
�N&����9�9�e_\�|� �bu.G63��i;4��������W�I���¢��̳�hw�s�Ny�j�^�;����X@R�̱+Vo\-�$�����:�ݻ�c�i���s�����Ih��yA޾��l�����J�U��P�@޶�c.ƺ\7�l~{Fgs�Cy��L�0l�p�:X2u@�Iohh��~�R�����e�i���/�M뗏
b� �A�X�#���P)�x{f=�\�[�����|J>s�a49JH���!HϰP�<������T�7��P�Jҁ���ba���I�z��2ΡP`���θ^{���pZ ύ�>7��5��m����됤�w�X\��Co�}8�G���_�]���M�XtC�#��T}�Fj�ϋ��L��#�棤��~n>� �7;�:�6�g�OO����>�ۭ�E䅹����wᄀy��6�]���q���o������X���.N����DvPub	����j=��V����k�4;h�jP�K#��}�D�VC@'�v-�ցd4*L�`�)E�J����}m	rYC^E-"���(!���U�)���n�l,܍���'���� Q���HeФA$��M�߬�C����R���G�ѩ 9x\x�{�.9���N�71��@e"��F�rŧ�����g`�,]�r�t�w�oHK� �$ `�k�x���iY!�S�7��%4Vn�?d뵎�K��8��MM1@�)�sL
[b�Q3�v|��?����.G�o~$�3��KN���kpPe��;w/���=��A��o������W�䱫o���+����(7Kd��j�I����>��}���Ƿ|�t����չ�d�X���V����&����I�I,2U�P�� ����$��ELz�i%�0��X�fSQ vI'5�Y���=7��A�3gϖ�V��e�$ 7�	*��zo��J�'���:�������F��S���XU��h]Ȭ�qt���w�|��HuO��3����5��=���Z��䈆�&=J@V7�ݿ<�i4?�mw8!�nF���={@����⚥��l�\@�m#w8�6����'�Dtm\5��O��B�o���ޘ&���WVnѾ��z��5�9��^NVVV!9��g(Es#�/�{]��n���CR��d����{nL�i����&����Hh��d_Q���?���ԫ�?��Pw:�����uK����jP#K��W��.��AQ�Nri,�s@w勍�$�����nw8���g�����N���4��A��o�e�ՙأ,yx�?��|j������3٫��sY$i�{ߛDXC��s���]a�3��˾�,Ve��Q^aII	IAc£��$V��&L�9����1:vP��_�������dV��`4��s'/i�PV�8UEK���1��Ns�ǹ0��fᄨ�}O��T�(����u�پ�zԏ���� ��]����>����w���]����v˥}��4TU�6����k�G�h|���\!�.5{*~ �FM�̥�D���з��/���U�f��"cy�2ٶPB��ѧyw����i��h�7���e_o��}�h5o��T��QUU�M���^��C���S��=$uh��:+�L�����[�ϡW�ج%䔿Q�w��$}�T~ k�b�o����ۛ�����/dp�x4��-�x"��ΔZ쾹�����Q�cO�������~=d�L��#MIu�s��Vwǧ,Op����o�����w�n���;�أ#^S���Z�����(����)1#^"l�[��M�F��@���r���:�ֶ�)�E 9�!�L�2�(���3�%h�#:U��}�uzvEN��m�34�r�v�Uh��]4wi��@6������޶�*�7�\�BÖ�%��!:=ZMc��EV+��[��a^�q��g�f���MM?�&"�C�7�Bj���j�;���V���F��	v��TNW{s�G�)-�m�wM���j�1��W]}s})�i"7�1��P��m�]qiO���\n7�D�I��P.�E޾=T��O��=��1쒎C�d�zh,uL��X(�3Չ>��4X�t<"��u"@n�9=؞C44���K�R��Wsۊ��XKصF8�{ʏ�rU5�ęKػn>J�͜J�d i�򼨨�?�HZ@d8�)%I��H�.�~#y���EߒY4>��??�U��u�X�k�_�%EӺ�R30C���<-���@����f��a~��'%�!��|�uӣ�cCH+xo���<�i��dv�xŽ��x�̊ə�x�n��U��HF�s,찠.J�pXO�m���N�&9!�H�|��@�L���&�c���*�y���6E�H5�M�KzP�3�1om��o��RT �R�O��Mо�d�2:�tF��DF�e(��v�p��B��y��D沷�ޔB� D�ㄅcZ1��vf��U�(��q��T�Hd$�}�����"������R�Y�T��A�m6���JE�OloM4VMT�qS��n�ɰ�,�i�ߪz�gs�N[�n-�o�$h ڸ��Z��q8�w5z��~?L#<�r���y�1�Zj�:j����aXDДo�5�ξ�B�(�ARh�E��y+&��kC�~a��l�
�����z�eZ�=f�s3t!�0(8c���PK�4Pq��W+��D���O�|�E�tT9���s��Ӭ���*}0t�%�M��]=m	~K;��?���"1���W=~��K%W�MN�m�r�w�$̐3%���9��K�����`�3��śWu9�zR��q�����rL�ޥ���f��5?������r6���t��Wq��PF���l������()������M��@��?i���bG��ry_𞊾�c8>�i��w\^4el��H�ē�?����4M�0Hʛ��K��eC#c�m}�e����O�?��Q�d�rL$�Yqd���B��WO�	��2�H�x&?������n1�R5�N%��q	h*����0��U�<m�N��G��`��$��"�f.ew�`.5p��L�[�F�]`V�#��2��AƷ�b�h��Y�����|���~7��VХt?W�4ʑX���F�4�y��|8[������Z�EOB��ڄ3����i��ʦ��'/�i�:�����W���Q��7�j�$�_��
P"�kU������7����.���ؿ�x��%��z5,l�%���;֔2v��h_MQ����N׿�A.������X�I]�88:,�%[�u5=XK��)���Mc<Du���YY~��"�X)DH�P����ӷ6>��MM[�����%����I�bI#��:)hP���?�"���R:�$��8P�ZZx,t�1{}���e�Ȯ���Z��0����S�����W&J �����(	vg*Vj�����%tӬ-����<�yˤ��ĝ�I�5]��~�;3���^�]�2hR���#�H��{s���lU��|vL�ۭ�����!ʒ#��d&���W��z��o4-� AOު�:��.��>��m��,����hg��`�@�>>e>H2ν�a4�J�}%/a+-�W���+W�Y|{���k^�MN��#�I�e"W���">���ۯ�;<��A�inT���]�0ɕ�pB4�k�[s�9п�)�.VɊӘL�}���0r����҂���qPn��{5�Z��W��9ŵ�i����!����08�x�r� oh<�JS��Nٞ��P�ZYͣ%%����UN6���������%�W��*e51�2@=�#F�?�/���*�������;Yŋ$�O׆6u��'�r���� Y:R0��!%���uV/�{��?<n$�α`���/�nTHbRA~�v\�ĩ����b�1�����a�,�r�S�������@�a�n��>R�X4mL����%
9�|�'_!����q=��n�ii@��Og}�u�ܵa��\��$�ߓ�t�N��ۭ�a*����#��͟�1htub�C-e�A�.�M�����"Er|���䈕��s�zHO+D�-�n��
��KP@V�c�[�ciE[w6}��r���{.7����W�v+#?���H�ʪ1��i�~mx�_���箲$՗�U�7tbN1�b��b�IN����i��hz��M��Ol�͐�QL���%�f̨aݍ�(��ңX-�5���9�<��ʧ�����:�Q�jE��쾚��#T�սi�&E�庣:�b��c�5����h���#�u�|�@s�*K�c2&_���!ᲁv�2�=�k�)�]f��(�&�X�DV&���ѡ�Z��N��d�P�v�I��w�̔4]Z�I:0\���ԉ��>�O�cЅ�[��X&Z��ۜg��FN.��d#\�����6r�[�8�j�(�������8Į����{���C����>$QaRx�m��/Lja�c���ND�s��,�q\N�5	�ެ�!N���1SL��蓳h�F#M3�����H)�>1�>eX�CF��R��\�"�^��1��7r�5��W�-?[���Z2�75,��k�ԟ<��	�s��d����
@����LV盎j �SX^��F��q�R��
�L�ҏ�OؠP��Z�Y������dc��o��.�>��Z*gш��C%�fn�U�T���S�Y�Q�fބhE�JA7�!���eK{I���6��uu1x�u���u���ӗ��ik�dV��>���,��@W����l<����Կ���c�qu����8�;�g��7����56Rc�r�d��1�	����缾�'���VA�7�Qޜd|�X���W3�)�b�n�7�x�I󔦐>�U����.ᬧ>����t���* �A��>��O�w)��6�Nx�_^[R�n=r�&�拌��P�~Iě/w��oUe�Hj��w4��t�GV��M���ڥm����ZD
,�_R P��8�����<����@��q h&Qi���T!tt���ɜ���o(	l()`�[����e
ce507����h'��� ��;0r��ܨ�C00��0��K��R8+,p��K�"�{ճ=�#/SN�]5"��_�ʏ"�n *Lqy;����]��kGn%����ܼ7���ߴ�0���w�_��*S�W��D�=|�Rf'����ܙ�J7�*���}��m�@ֿ�c�<5�6��	���� �c����+f���	���%��Z�fϟa�}�9F�1XpJ|I=�Xk� �����2.�W�_���∧��eei��v���蒘V�Y�=zϟB��/���ډ����ʗ�Sc
���ݤ����}���.A��|<�2�����/��h�C�z-�!y�$��Y���3���*�/�u_�N��ߟc�85��Ss<Բ������������i[�`���?~��1�c���������_����NK�Y��(�=�Ufu��_ѱ�1ã��m��"��)��kc�������'��[v�:�seד_o7���7}��N����WI�����n��V��A��;E�7S�7���>i)ر-�0��<!�c�������Ҟ�����C4�$s�3�;B%�K�ߪ����n��C^-]]]��B.�ub��/���ա[?��j.l��O�&V�q�Ӧ�7�t�������N�?-��y���*�Ґ)RK��N3������"#3L�q*�m���K�ܷ�
�|B��~!!܈������
x��R��֡/��4,k�$�m��%�t�;�u�U���@۹&���neWA9,�peP�'`��R;*��ۣ�>@�b�n��,��G�v�;��p9#SՒ�?�BVr[��D51;��4�]5E�?�������������S:b������'�[�ޘe��g�������q�Dq3"����V#F��cD��yS���\{!���ia�"'.'���A�A�`���&�+���#Ԯ ]Q�^�X�"��j��Ƞ����i�e]�s�γ\�?��vy;-�]�cB�g46JL��n5_B��Ď1�[,f�Q;��D�76�\���2b�p'�s��/&�90b�p]�.F�U��I��c-��2Q�-��}�����0[G-.�����0�%qc��/x�B8���it����t{�Zz<�օ��3�[r��)�z`;��Ґ��kW�r�>}�Qn�H	��7�����SM_8�hh���b�K$o��)��y�Q�ccc _S���f���5�-�'�o���Hi��2�� �|��K:���~��������9��t�����ᮮd�HΔ4߷�i+����G�zF���'x�ϟ?���� ���u�ze�"""�4C��n����f�i�JN{�ol����-H6��cuttT*;�s�	_���`��vvu�;�h�%Z�K��7�av�n�b�
��mHC��$][;;.ֺP�.�
v_�mvvv�@ �أ�H��^7;�}3�_~'�өkok��(++Kxt�p�r%���>?,��hJH������`���������~~t!;�~�"�]N���9#r�a'
�P���-���>��{DF�|���"�=ʭ����U����~�ڡ]���ګW�����+p�w����(�{���\�.��`����ʙ[�� �Q��ի�(N|�D	�PҦ����}�{
�� immm��B$E�P {�<_����|G �g���SIF}�5WG����#y��X�!8���Ɏ�;�� �ؖ[���|���-0_��,��{*)z��� #�EB�qq���t[��s�u�d�m(�[s�s�a�c�s�y�8�g2��t�����1��雂����y�����3J���'�p�B��a���GG(�5��8�,������Ȑ��~�(��x���*���X��8k��b�b�a#1��T���\��[�T�hn�qz�E��NL2�V]h �/>-�E��m�2+p�U�tڝ�ƀ�g�B!��>�&���z�Nt�ꊭ��j�p���vm�� Ij�fu�T`��e%%�L:D�;��n��E�/���[�
1!$$+<Kj'�⫺���Ъs�9�`t+�w�V�#`5�L{s����s�#�D��J�B+%��)t�3��^����ط�̓yQG�*r?�	��~Ɍ���	ؕ{�m��?~��Bd�����Qo∓\Gi+��>��*���P��h�dv4��b��b�brX���5�2?����
�����d��x��Q��=��
JJ������c~���Z���(��z!i��������SRRr�k�g��@"/�z/��eqq1qL$X�d~󼶶d1���gVWW��G��F���.FG�g�������7���l����d��M��a�kkks�;J�j�Վ*aA���/W���p.r�7���=�9ٕ�pػ�K��]���~|����|ž{K"��^$ykQ#k���2oƢB�ŝ�Z4e���4���s�̓;6o��ڵ��V���,��z�"Z:ƔnQiq��h�< ڄ��7T���}���ǃ��ip���y�%E�B�5�6��F�[t&Z�^�l<3��|ƺ�m�U�:554E�����O�xَғ�2�i&������A?&��>j Swv-��|���`&h)�3�6��^4OL����i�2�d�z�~v�$gYk��*tU�1��Gq'��;p���V�M���,�T�x�{�
�����+�m�
\���0�K���7ȎS�Q~��w���=g�{�-z�n�3Z>�g8ߊX�w�C�z�͈Xy�&psn7P{ �
�ʭ==��a�s��LLZ���4���d_w�d>��JV��>mU��6+e�i�����C���%8��������,�(!�j���5��'�B�oU[?���Z<Ho���M&'��r���K���d��}���܃۔=\\N�E���cc����Q�W[�}���䭄�����#666��� �+�=���j�]�ַ)�q~~����h�I��m�؞t�oce��ȍ֜m����&�k��ZYZ:������b�?&�l�i�<�]Z���
]wBsA)|?@��u�P��*?�"��˃��օ-)>�GA�vYc������}+ �sI�G���br�Yy���Ѽ��H����~�S:[{C�ä�����t�\\\�>�(\e-�RX9	,(>W��fB��~���a�A}dU���Z�;`���Y�;��H�6�x����Y�h��� ��^nM�o���"����*9��͚��Q}�ϟ/�#�}����(�D �M}s;�DjC��w>����{�)%���
EEEE4�%>�� �5�{Mu��H*�W�M���4>V�E~�ۀL���P�\E�f���HlaaaO�@L&�2�p������I ^���w����Po[���@>�����{Ok��O�~u�Syg�m�%�)E(Bgd����x�`�8�l��w�7���k��(J����fI]�HP�]�N0��ĤV����hS���)��(�ۯWB/�޴����"~�}��"c����Δ���1��>CCC:D)~�ׁ������9��b,�z ���6nG*��(��/�)���Uc
��q}|�koҞӧO�}�%}p}(sm�bS��<6f_:��V�p���N^
X[ ��O������Q�	��
ŏ�qát+**��u�7v�3<TS����so^�őӼ��`�}�{��~�u���;0�1�QL�#���-�	E��$$$~�P�H8RPIOߖ:�ܦ�Mļ��={�duA�9 ����20��\[��ˆb���z� m���DDE�ʀ��Fk����3�Ү�}b�1&9�7w\z��/,��d|?l�������^P�H8��GO�ӯ;gs�寫G�_zg/��������>ם�C�?�^��zW���n{x��] ���p��N<>�[��r�0oOF���r�Z�\b"�&%�h#�i�c���~#R���[%R ag�y?���+�肰p��V�K
p���M���sv@ZN��y#�B;��/I��\S�7=�2�o�=�.���<�}���Iδ/N�&�9Lv?�YZ@�����ϐ���q��cԥG�{O�)dR�?A60��y˂H�������{��wm�N���ܑ��֦��\bt��U=�a�p��O��ևN��W�\ ���e���l��:D�K���{�ᥩb�g`D�58���h��4�S��	)<v��5G��|GBJ*�������n`��Pf��^d�.�l�MV����{�Q޽����t?B�s��a�6�8��oUl� |d7����[�*������t1�������2@�?Q��a!X*��;y�-0�m	( ��z�o0�F���5x���j�X����d�7r/�F9ݷ��WrAͽ=��g��J�·�/�6sŖ��%v�	�5wՔ���^�IS;�$��N��UUP����Ӏ"����K��K�2��Jan�o�;ب���0\*~F9����?�q���+���៯�9����.��J��h;L�dd�*XE��'-�^`[�2����+O���>�x��S1sZ{���v��<9�GƑA��k���96R��Ff=U��W�$8b����H:�2����?0u�5' ���z͓�?v���lz�u}�x��հt�]e���:�d���̓-g��Ո��߿vv�m�C�:�K]j�N�ɞ[n_��FWiw�_����z��*���m]h���Z��gT!����}}�D�_b�����e�cE.�W\�f;�?���$B�#-�=����~=~?���WO�>�sX_�E#)�F�-X�yDnu��ݹ1g7����	F���'�k�#g}MUHH0P��qK����,��K�a��r���OV��1#h\�e�Ù,�����,��A�,p
���"�M�; NJ�^�O;�l	���X��hm�SHHe�Sj9��׫�^�{Ⱦ�!���۳$�E�u�2P�R:g��A-�K�������#q��5�����x�N��EV��9Ǽ��~�;�lw1((�|�b��!��F Dmk�����e7���Tt����-ժr �f]�oo��J���3���P#(%�����8%rų�z�бN�^��[��i>x�l������H�p�u�(ԑ��������l��l˻�KL^	�
֙	���^���t��A	��;4H���4��ț��v̍��	�Jy�G}9��>�4�%�>g���ǭOFӃk�>�� ;O}}7��N�߿�e҃bF��T�����+�S�����<����yR���\A�(��T۞{l6��xk�ܐ�ԺY����y/(dM'���������z�-����j��u�������P�����9 �M���}��%�PAѻ,�H��O�qN3����id�*���6�L�8���t���dW��'�{U�}�2�,qhH~��#�� �gk��Kkkm�� s{w�uJ��4wy�w�Q���;�4<l=�̠5��/����P�.6�M��u�(�.��)m��#W�AiE3+3��VN�Nm|l��okkk%E�������}Ϭ�l5���&�c�k��z���dA��"d|窉IzM�w+�ɼ��g�����f�- ����
�Bڎ���Pj�����Ǐm���s�C���$VO1+N6����E�ZM,s� b�OyS�� c9��	�Z��ŠA�CEތy���SH�7	p~���[��)q�)�R�K�@��(��sUS:KP[]�������IO�ZAC6y
4�\Z_/Uh�/x�ж6�J�����@��*�cx�򱶒#��,Ō�������h����o��Q�z�5׆�*��o@���9�O�B�G]��T���g�$�99���  �y�e[m�����H�T\����	�-�R ���� ��f~�l�fׇ���@�P��@����΅�iu��x��^?����i7�s��FC���>7����UHv��&L���� ��Z�v��e��.���_޹s�]�������]�0����XѢ��D��������4DiA7���0�@<�e�H��[YXCܽ����6���LTT��I��2Ps����5��!}�&Z 0΋Ł���EAkf���,`J��Gj�<s�
���׽{�+++ڢՖ A��[�����փ𝝝�K"�E ѿFD�@�V��꽔Z�������p��)�G�?73�~�����\#����ct�qqq��@O�@: ?M+���<�E0�\��/;��ŏ1۹G�(�e���:ۮ�0ُee��Jjj�Y�_8�Vd��ew{�����b������P�}�#�J�����"�uا[�8���khr�C4B�*�l
m�LG�Sdd=}�y��M`���D��N��'oZ[G�'x I4@@f�O��B�5�{���E ��>*A�&�� ��`U��t�КNL�Y\Z��R��Muuu�Q��� ����
����(3Ͻ�z )�<w������9y��AS@��3�RYV���np�^-�j�rè�"1�aE]�p��c�@J)	�1<\XB���K�@F�G��~����3Y�q� ��R�;
@�V�� �F�q�8�5�M-�ǛR�]�u�H���$��0�z�|�f�we@p�PD����p4�Ȏ�3���5�Y,0O�:�� � �W�]>`Z��u��; �W���<X~��ٸ��l���v{v����#�f��]0X���3���t�Cj�^(z
�k��ʱ�#�:��,�l�w&S�޼�����>��Ό/��P��Lɹ�ӿG��"��x(x���=�/��U凈"~��!⇈"~��!⇈"�+�w�Q!Xz����б�aOF˸�	��K3��qTMi��2����}:�k醁١n�r�p%��k�B�{��r�\W�ź�ݺz"���*R'u�H�a�`����
��Y��\j�K����Rf(���(�>/�7@A�C�~���������X)��=���pE	I�s�x�@q��&�pbS�W�UUh"���XcsC�,�8!���Ե��n��"�}]����Թ��nj0��k�>����$��U������b������XN��Iǵ�P��Fde��]6~�������챱t2b�"��dG�������`��nnmH�~m���b"�E�>`�ѺЭ��/4�����(�7a�[~@�N�2�z)P���#\*����]es�jj��E`�切Z��Ue&��y2:H7�qgȄ鉄*`	��v�C�ڜ!/���c7�w�%�k� u��%''��Z�O�s�!X�����.�Vc�XY��쉿��^���c�;:�k/>0$�������dY�4`��>bG��V�xgw}=n�Ψ��s�N�����
_����Ę���Z�?(o��v�Z����P��N�s���;�Q��kG#Wm�����C�>]V��>6���!%$%���Y�U�<.[]]�&���9��#�n�+f���g�O0om��<���(�G"�������PK��ƚ�Y~�����5U�C�!p���y�Y+�z��rO��?Ǹ�`=~��~^�Τ�54�ھ�ޕ� �1.e�KQ?-�3Of�J3�2^k�<�be*�<\kl�b"���xW谉E#�����Q�!�`���;W�l}�
��U~�l�y�v��W6�N<���\B�\^���jxH_�g�Nx�A�M�ov��"��Z��n2'�K[ �0��0����7&�ASH�q���@c�\	���@��h0èв�+c��!2{���L�򺡡ap���Bˀg�>��Gg�x](p�;��櫼��{i��Z(&�S}�K�X=�fCt�lH�]�;�&9*)���g��ŭ��
�y��˄���lxRp-u�OՔ��X��(0�m����YEEE��)j���)��A��$�c�=�tȋI��8�/,�8��ϾyWZ��C�����-""<
��Z��]ʎfu��aP6�G�,6ɒRV+ƒk�Y���/�
�� ���t*��������DKc����)Q���4��bͷϬ3� ��i& ���!�N---��T�"�}�]��k�֊�k�B�
��L�H3	Y�!͡��.�$��]��9�d�k�f��jQ\+	��z3b$!!a}�>eN���ۯb���1��]��� #�.$$t�+p-B�H� ��n��KN97bc�80���=Պ��H������V`���#8�~��Z�ǫ���-#�`��ަq�[��2R3,(%��⁀��0�«�.���)u-��ȴ�@1+++:^�ߔ��p����̑&��_h�-d��Sˋ._�$P�k����E��m&�@Š�_��ɻ���:�HQ�����hR��NJ����Y�fbM�hȫhf����G[ر��~ZM���!�	WBta��FG1�]�U�chh�Ҕؿ��]3	ŗy ���\{xh�M�@�d�;�A�ݠ��f��턃�ە�FFG�|�E��������8��w?�`�OIa/6�,� ���3P�����[�o=i�����{3�]����m�ģr�p���6 �6����I�;��h��ǖ�!�}�� M����~9�-hHs�3����u�t�0S�9����������n�C���D+>e���� ��6���QÛ����hZfi٦�`�s
~d����Q�7�/4�=�P*�6�_�x9�{>����0
��qg��)�v}�yZE�cP���NP|�y�Ɖ3���a�}�@&gyY��dX�e�(`~{��GKK�]�Y�ϝ��\	�{Uc��v�����h80"�7h�}Ҩv4�cA�c?Ԝ@�
0�J27[���'�]K
^�i-���� @F�������P8'�Ӡ�s#�u�Wjԣ�h����Ug�L��;�H��P��Yd��G�Nr8Y������{J!��E�fKl��Y��WYg���@��k�9+[ ��a��½1g.%����=��
�f	�w�N.K 
���`�?�U�ܺ��B�m��+�(�Cg d ,�s�
z8�IZ��ʟ�jqZ����_���g�f�l:' PQ�NL�/w��9�͐�� ��=+tM8X�=Ҷu���)|HK�f���<`p'�}�.J��<�C*���S ���\/������7���d;�!H5%�+S�]�n&�1c����e��K1{ (�[]_����w:��Wش��������q6x��U:u�DB[e��J�s��a�[�="����W]T*N�حK;�x��H9'���`5W���)����[��B��.aU�h���rz{b܏��l�����w?��p�Y�Lky��@���j%����W�h���_`N����ኗ;`��>��K�{Yh�3G��A��.����x[�Cᑁ�/2z�p��!G�c��s�-�"(܈�ozRK|-<�j+�t���g��E6��5�f����y*��p%��}�7@��6w�~ٻ�����m�ޅC�����L\�y^,��r~���q�~7`�"�#{Ͼ�0�t�&�}C/�y�5G}�9� ���I�/H�_��� ��>�tj^�Li��Ȳ�J$��"��.�l��|�w��iY����妁]�8��0��x��)��Y� _�?CUuu�� 3%�V�xpk/}s�B���l��p�������I��3q��AP�n:�*Z����
�Z�OMKK�i)Z���ˤWNiLz&�w-����H��BK�!@2�~��Ď�� �M| wwG��s:��Tu�A�-������H)>+�'����yH��d9;26�"�k������h���}��C�W{��d��Ʈ��`C��8J��#E�2�� ��&�Gqi����D��&5BD�R���� !��y^fͺ�Z�s�|�����<��ߦ3�O�3L��^�����hhZ�z�6Vb�[� �p���]�1��K��>��5�
)�6���r�0�o��yd����p�n�� H�X�N�V��zV�J�N��l��$M�������D�Y� �3��U ٤�3��x&U��M�I��x�o�}Qj�,Jg?'�o�M��^`D�{9���´�C��'���v����0l�߃��y���" �el�<5��`���i�zOT�$�$�MX�@[D����S�Sr�D"C�3��^��� _	��?=B�ӳcL߸W$�W#�cr�n�)�=BO����|�,�$0��2;M�b�%C�h�&��ts!��]�Nۃ�oq���;�T���nXl'Rގ�{���3m�����>��6��(��^�)�~�O�'���y�z����g������V$�ާ���^���񔘞���{0,�kV��Bqɴ~1�G8$5�OF�A�s�j�C󙮅�Ӣ"��.*R��#.A��j{>�20v5I+*��g`���
��E%Ro���g��^b���M&�BR\� :��Yg��B�y=hʸ�j���=Byw-&l�$�(��I2�`Y��Wo���k���5Bۗ� o�cǺ��3���K�t�������`8EJ�(�/E���nݰ(4-aF�5����:D�?
TM$�z�-��%Dbz	Cڀ8��Vo����X���*�Ͽw�#��hƊF��N�d��$\R��oDKՖA��~������ ��B���uW��ާ�N�fԳ�7�<vD����"�Qg�x���M���ȝ�X���u���:��i^^�;��Ř���w�����Ey�kⵘ�j��z��D���a�y�ު:_Ğ|_�o��6n��j���������8�:s���DW֧���X��Ƕ���N��g�.�0;H�2����Sń1�U�'&�����%U�qO�g������A� �3`�^5;�����ɋ�*+�zJzz�E�"��@S�4Pv�/�P�2���W�������ʾ�W�L�*@�'������������y��& 999�e�<�<��F�W��s5!MO�'���co�t+��=��o���b�̒��gi�/�H*�&��UU���RI��3u<[�>�cVN�µ2���|�1��ƸsVz's����h`��K&��Gu���{����&%3��^d��Ui^����L\X�r.�	��{����|��Lf�h?pKm�ڳ��NW����s���{��e����[½�abjiam��s�vT�v$��2_�k��k�K'��y{��ڢ�c9#A�E��a���yw�2o�Ac����NI���H�7����q.��qN��Y�K�����櫸��i� dQ��&,���j����pj�gj��5#��%ꏿ>�d��R�r�i���s�*F*U'��$�"�#�H\�F�i�F�07p�ټaZ�7�o�����
��R����Հ�~��#N�vH�im7�VR���6��{�-�h�#�T&�vŔ���19}�v�O*|c,���{�Cr~���A��(����9��eu:~�:Τ���J����~}\��)��بw�eMƴ�4ѓg�D��|3 y�<����!
>I�)��Z�uXd�>�<�|U�>��b�7�%(��q�����m���[���9����k�bы�N�hu�o��3ms!ZK��[�M	�n��7Ug�"S�ݬKfe�.�;�;y�� �W^�^��]��p*`���G���(�5�5��h�pss�n����p�]2	������K�:�վ4�rE�̄C���i?���(����90���
;�Z--��Enݠ�
'B��Cǿ}�u�<���������;Z��8Z�*���J�^�xy���a޻�4�Fp*i��1�^�W�׶����_��$�� ����)P.�|"�"4C0S�Q��5�;�ױ�b>�ߙL_ss��_��%��uR���l?������>��mm��_{��h�^�dg���C��ڴ�fa�B3OO�cCC�ݾT,����[���%lQ=  I[�Z>pr���:�`�R��ه�����J1&���|�7O�-P���������ԳV��!��IA^^Xɡ���O�|���I�����ź|�)��"��Aq��|/ɼM�8����A!R�zm9�G����g�B���2�ݻz�.5!��z�Ӳ�_���ܸԑ��o����X}}=�����111_�;�ۃ���kGy3V�c7X8p�3f]v��i� �oya�_qk��8��L&猦]�tJ�÷ډ�҅���oł-��͟e���ڠ�jK�f�������,��@�0[4
�,�y.q��p�Fo��jJ�&+�x��X�9饝��E�\h[ ^��oY>���*�����S��p����x /g�������I�Y\K��j5����۪�E=�O�2�0��f'�K��K���7v�� ����R������)���6 U:k/B ~�j+'Sٴ�jv��*()��ޝ/��ml�%�X�M"���F���7{�iU�p4�wGm�~v#Q���Z ��������H��5��j�6}�sc,���0X�j>�۞�QX�����������2l�D�rݢ����� �񂲼�$�M�0*3Ќ�Z��(tyC|�>���9x�츒����V�� c�#��vS���VG�Y#���0��s�z��vs�,3���G�⦫��w�0Ot�7Н�D�f{��A�/�q8����hKX�s��L@J렣��1O�uyBb b>:::�*�Q~��  F��irgHj� :((�|���@͊q�K�O@Jࣲ��ic q���u�;z��հb��#%�o ��JS�G��VZ
��U�1Ґ��	x�\��&���p
|���D����3�R�6��W�.�p8�⭗�pv�G�.E�&�7�Є��K!�󹃂%����mߑ�B�F�d������A��V^��d�2�O�5�z�kZ��y%_��?p)0��*���*�
[sH��>�q"��Y)ۑ�0����x䔕cT�7�0D\�q�	@|!�f��ģ��o�ۥ���p!�WJ&i���l\&͇�^�Q�5Fv[�*}��hPH�Df�D�Ô���7�O�����ֈ�]|��y��QZ�_u2��X���6]��RK<]�9�E����$'Զ���F��Ҋ^ڗr
,�oo:P|O��E�W�Ƃ���Lj{�K����j�m���8��Ed�F���o��w�}�r(��:�[La#`L��-�	�[[�����x��`��T�d�dh��N,_1�^����|�[�e��S�C�zY
�S;�{m��`ΐ{#���j��#9��&[�uy`�ᚠD���!�I~n�y�"g���e��"��Օǭ�W:�תjA��^u����yߡ���,���\��^���U��7:kx��'�*o�3�::������L,-I�0XG���k��w��qyJ�c�W���,��#���r@m�{y]w	����Xg�E;�S,^�v�#�;��***�c����WC��Â� ,#���V2��3t΍��Q:9ە=�='����>����MW6�̘��E����T�`����@Iȓ�Xb��ӗk��G#�(��S�v)CC�5�tT4@��d�"دrL�6�r
�7O��э��*�'?^q� ,=�(�\h�Cv-��;���5�H��%.�,�&#�E-���'�!3�4�=x�[ĵ��>��N�o.8�]l]^��h��=mPr���V�g،s9isac�g��慉�UJ!���Qh� �ޖ?nq�O�T�0�wyK�!YC'XB$�h��Y��#�G�?����=j���0��,C<��C����%��Kq��-H����!�Y�1Y�aU0�̦��z�R6;�,s]g�?�g�X�F�O����3�W?�GG䮃]^Is�&ȁB5�<��t�ر����ե�.}��s�?c����,�w17<�����^Y{�)��.#b^�����t�v�4��]djIN�LR�l��0�]�(���p�\]���
��U�jGp+[7=��J�rbT5%+��-O�a!F�*�=·C�&K��PZ1�T(g��7�.�%i o��jl�Cg�B��"߳2H����D��L����Q�k{0r]���6s�c�LG:cZ��DH'�K�O���~�}<�U��&���!<�����sya�'rV�p��'(�,�U7�/���TC����U��AP�R�Jxߊh����W@+u@MO1� �tE[���\��tga��QZF�� �*�Sh�
h������9$%99�7z�yg�|@ޱ�\\-��Կ�,M���C��W���
MI:��6�:�t9om^S�V�����Z�n���I�{N$���Uޠ��0*���!67��W�D<�dΚwH#So�*�����[	h��7��V�'y�5#�s�k��
m+���ǭ�^'��XY�+0m%�@P�s�w~Q�+�D�����VQT�jj��i�v�cÊC|�"� /N���2�U>�|�������X��]���̢.��2v�5gN����ا׊�?[�Z�Y�p�Hj������,t_�Pp�����`�
���������7�!��񄙎�������s�쭞Ʋ;���~Z�u��SZZ�Υ�z'ȃ�֤��)�U�n.�1��f��'(��=�Y+,���Aܼ�M���l^�]�uM^Y�|�c�[�������&Q���E����;�8��jDG����A�=���<z}�
�^�����}�;��֮���$���}����j>����Q������M�ϼ�س����I�ų�2nè"�`-�˝�+�J�����%��[�<�v6UL~�5I
�qO�����J8�31a#Œ��5<mx$��;T���R�uV����c����
����ŋ<�{1�gTxWd���kH���nh5NP��bɂQs�a��͋�_"fyQ�?@�#�c���]+��V��[li�VX�D@Փ���c������Vw�p+z���]�/:�ƌk���9+f����x��E�'�h���F�v��/a�����߭��G�c�d��g����:6AvL�����x5�/'��f�ȫ�A9�[dpd-k�ު�B���!�+�AJU"!����7�JF�Y�Ӹ�WKl�_�I�VH_O�b��w,A駱Vv�WR`N���mKeR,k�'-nm$��X!Tl�]Q\���%,�E�*�-��B}����辒��C�=�g�N� ��r��M�S 	:pڇhืE�p|]3�2��S���xM�h�� 咕��me�?�H��P��9
�n�%n��n�A���7��P`�,���y��Ϧ���b�`xdt�Q~C�ş�m<�yY[�+����Z�#3Jxlk�8�����>���%��Fs/�Tm�g�)�P��:��(�Q 3�,�l6�v��ds��&��{zQ�'w���}1��DTw���	��9_!DBߩ�TT.I:��]���m��n��Ǡ�㯵u�,���a~�4�����߬m��T�4 
����w���z#�m`���ޖ��>нUtx���������?n��ΒϿ �sb���ܧ��4] �c�-\�%��r���N<@�2�$_��P�_��I����94mr������|���u��B�.r�===�B�8o\�륲��9����������G��+�?尦 $[��a�ew�9QV	H�����������p[��� �`'׃�����45'�u+�S��Q�,^����0?��w��F_��a�(�G�,Na�SR��Po�A�k�ȶ���vz5����X<35u�Mv�o�sӸ��Pg�^��7�}��kBd���b��ʟ��ځ:��E7�����2�������I���݄㣹�>��96��T�˴3*4��R�����=���D)p-�E�u�,#��}@[ڱ����|wے�v��������^���b'e�r�p_���Z��C�t<	�U��ᘄF��O>�v'>r��Z�I�U�$V���=�h�~��٘?[��T���z>�����ѾC�dD�=�4v�;�TN�*�Obܻ�]��5{����8�C�5����`��Yk�,Q?�*������]�����S�I��� �g�U�Cގ�̃���G83�/#��^�ea��D�[��~�b>�ٗ���7)fZ��9�|P��F�+�"�Rt�����Y�iHBq��3b�\���y�U;I^���7���;��*A���w�e�oҷ'yd�~�%�.�r�P�������{��@#�S�f^�qL$��F����b�|98=%Z��冘��iv�kC�'i]�r��q�N��@�Y��tr[�K���Θn�����rk��@*�W�����W\��P�-Kyk��ӹo��ӏ�y�B��c�V|����O{WʶϢ�g�,���&fv+���ƭ�gBY��,z�_L6��֥�/ӝ�����Bt�`\���M'�IcI�ǯ!�ь��&�+rs�&�λ"n�>h���]�j�6�IOrzzz�MԏS�'5QK��Bi͹,p���r(y�< ?a��t�L���<u�y��*vicѱ�~}�΢M>*<.P�Y��T�C>���4tS�ڮ�H�0�襁��lh�D�b�^yۜi�k�v��NUYV�k
E~�/�c.^�ҍ��c�<u��D�n�0�fI0	1�־�T���X��bc�&�o㳲Fߝ�'��&�Ag�(��kf�#,@�`)�g�q�lfg�w�}ou���$z:��=mꂜ�s��N�H���n(o��K-�>�]`d+�,z[���4���N8Y8z�E�I��|F�w7�~ȹ��� ɃS��J`�Y�Uz�hCç�W�n�6�D=?#(tHi%���&s	H�w��͋c�{����<T�(W��qT �'}K�R���ҳ3z�qM��{�C���]3�`�L)������Lp%�;g��֤m����K^�3�x���}����蘫`o�h�_k�f�P�U��m/(��a�*���4��7u1@� �����f`�(�pN�3bZ�W��R�:��du��/�����%O	*���؃B�j{N+7o��}�����6���a��S�I�"���wuu��0)���8����<=�5�Lf�n��TU�PV"n�\��T77�{�`�_{��6Ԡ�h�L�	5�|��{����ג��]��]�J�������]'� SxʔRuMY9��(���LB��L	��Y�������(���2����r�\^c�W $|A�P�/����ё�¶�^���&��
ζbt��$N���|_I�kJJ���3�青~��Á5ÑŒ9�S�Y2b
�:p�ߺ���c�C�S �>��x@�
��l��,H��
Z��Uinj�e�LUv�����������:�串@�h�So�֥c8�������R�),��R-s�1�E^�P��OUx�����6�ɛ��L�ο�T�Z���"�M\�܃�?�X���^F�.��[��n�k�y��8:D��������t��>fdڞ�����V/�뙹��)���~��_���|� ���Qqk<�� c��U�d�Dp�3����� �:�|�
d���c� �7���-�����kԊ��/�2t,�����x���#��!�R7�U�|�^~��\wԳ�2������,L~�jwV� �3A���aJ��վa�n�;�v'|�hGؗP�)̻����U���?�T�Ay~O#]�P���\�/Qڜ��� i��>������������:�}`{��j��u����Y2I��1&�4��X	brʂ�-�lv�;�R*7S�%o<��_QQ!2�y����w�������E"L���dKP��3G43;����?�Xy�4sO3�K�H<��\�%XY"�s4��| >����Bc0�G��%�>��Ny d&�0��g�ų��'ےe�2A�C��)�j�=�H�����$'�������ǭl��Jׅ �b0&an2�fnV�\���q�q���6�k���{P�V�hsݗ�-y܊1�-�U�@H �%�f�2a�30$��6$�;t�W�
���S����8��~��O�<M��1���6����*��ϊ�������;�f[�����I�����3kY��d����g�SP�tu��MXyՕ�K��n��=Χ�̯���C}�;>�i|a3V祡�an��������+���:�����X/2�?o�[[]��d�t����ͮ2d�Q�ם��n�B���/���444��O�Q_�|to�����Z��7Pd�)����I9G[ڦ�mp*^�������,�Sٮ�OYB�����a���?fV6 ľ/�0\��fd=0m�[,ȧܗ|�K�V`|�}XKmN�p��j9��*��G{�a��/9��9Ŝ�rԨ�B�f�
�=ٴ����g��΢`[߱�<Ga� �E��_<�6�;CB֗�<n����޻�^�pfbi���18�˅9mY.��[�'�H_����D��7���h��\���f4u���y[��H�B�rV&�Â��M]+�y{��W�OY��>���+�y�������W7���1�&cW���lYM�1����g7�O�<j����A*]��&�r��2Q��̜�Թ�0�����4BO������.��6+�-;+����*�Y���](9�
�7,H����=��r7��@N3�N�����w)�b�)皇t�[�\4�f=HmK�?�Ҋ3)0*~��ߺ5:z���5��}�J��I���	��2�n5�L;�	�^
��up.�"6a�(��7��Kr�B:�wH���onn�g^�ݽ��KD�P���ȭ�7!O 4�Tp��,f�^�<R.E����_��I ;���Uij��3(.�em	Q��o�+ S�gIY��r��x�R.َJ؅�� -�~�O9���[J�֥�|� ���l
VV�3ȝ)V��]\����1g�3K�
)�;H�H�>J Z�$W�X�R|]� �?W@��Wi	|wLO���#���W�5���MF�$ol�cȹT��#���N�<��x� ��,CC��v����O�q�g�6xuR����(]�zve�Q����ߐS�Ǯ{Ng#A��`���Piq�n�\,V�:P
����:B�m%�a���M�Us�ﲛѯ�V��2_�|�����I� 'O�����o��	�P�G��y?��ؙ���\�`@�iC�ű�Ǡ��N��R��Z�C�-kxz{�#:��G�g�륹}-��-�k�%_eu��;g��g�q3Ο��[99�B��>u�#!�ɇBa���� ��� ����xX��a�!�n1��U��������h�_��Z3�Kj���9�B&�:�aꑞ��(��Rb"ʶ�r�t��xiJ��R5ަ#v4��S$�;8��đX7��P����F�op��/2�P��{�h�Nz�^����0p�1�E���m����b����XB�v�{I�ԗ��7��4WB��/��^�v�N6㵆�U���f,�0��'[Jf@AY�Z-�4�LSgC��W�>�]#z$f]lƀF\ӷ��o2=�z���q@%h����;�9S���q�.R4ֵ�����)�O�L� >9�/紬�W )R`DY��$Gr�зJ��D�ٻ�ރ��*j�V`*��t-,H@���+�g��=�e+G�<~����~铩���֦�T��P��{���@��Z��e7n'�䑐������C�8�$'f'C�ݾ!kz�=���T���,���X� ��qOv�튝��ع��}a�����m`����9�Q�G�~�����U�/�/�h���>�(���?
�(�t�ط��(;	��B~�Q�G�~�Q ~m���Bz�����>�ݑ���N����~��̺��&�p�޷{�9�=����=�ws~ϻ�ZpA�M��s���u������u-�,y���B��i�g��OM��k#!s����=���>(�G?��Q���*Z�y�W2r����G�R�������2��B������ �]A��/s1V\�G�6C�洐�V��<��kV0Ο���ءѾ����%�����VQ�J�?��0�0��%-��7�=�le���k-�3�5+�F�SSS�'P�clP����X��A+���V�σ�G��ʬK}�>}s�+�8ʒ��~�mh��Aݭ�ݨC���[����U<�e1�}_`�B`Yo�Y��J���޿X�� UX9f��F�.ߒ�W����y�+�Z�e�#d���Ӛ)�h}�����	�%�%Z�sXa�w-y����Y�X^�V��w��h�����?����Fө�L���K�3mK�f3)�3�|�iy6�q��TMx8�2�>M޿�\��P�d�#̏�T���]���+�L�v����tE����+h�z(!�wϢTg!Cw�^�<[3,"���P�8!�5���*�Dk����	e�\�9F���#]9d]��Q�Ec�Ț"����k�h�Zq��i�򲰪���3����+<*�����N4hTj�|%�� ��F� �c�]�x ��;4˷�]�k@����m��;=��Ѳ�V�Ñ�q3v�wp����x;h�;��|x�S��sPzX6Bu!4"�M�Ǖ#����2���5�WL����@^��:V�鈼��22<�����	)�:?6��~��y�v}����tm��ׯ�;���)�ߵ�K����"O�{W\̞(a���':xR���36�Ez��7�s�Y���ǭ��O�)��6��3�u�<v�*9��Ɏ3�Bo$"� �553�kii�MUX�(�@��r�"����cj�Cml2ɹס�"���D�����	nך}�s�<H��="����c_�re���!�q��nؠCW�yu#V\L����E�������;dr�������F�҈�s�
&c�#t����0�s乚����,��'���gT��V':���*,��+���#��7��aDg8�*o���H��Ǟ�O>+�m��� ��G�IOTCks��Ή[����M>��m$��P�hM8���	:Ϗ���wp]�r!68 ��O�!���D(����ݬ�NY��(�݅rM����x������I�CQ���v+N��@JJ*]$+X�_���fu`�Z��v�R�t�� �����.�NF����C�L���R�F g{�*��tT�Y=�_PK   o�X���Es ?{ /   images/58ea960f-8973-48e4-ae29-a018cd448a26.png�eW\A�.L ���-�������� �www��a��>Ϲ���8k�f�ݳvuw]Uuuuu�7y	$x|x$)IQ%��<�����o�]J�>8)ICTL�?|4�����Ex6���� �������0h_l�V(%*��w��}w�c�	f��=γ~z*�'��)Ę+�R1�A���f������l��R���
�4y��%���h������ܜ�`���]�O4�3��m�~���W%|2��-&���WԏB�s)�m����ϕWAF#��? }���ok�����j�*���VR|H6����4j\|�[�B�G��U�����MF��D�?���DK�rTK�/�����=���SSB�FO��t�1�	����"��Lv5�5P�ȞG(�T��ӕⰨ!��ˑ�{j	ؠ�����o�Ԍ�V+���5�Hק�ؐ4�o4Dp��X{{5��;	�	��Xkw̜9^�f>�Փ~�+!=ˍ=7����k��>���˷t|e5*8��l�/kϤ�䎈Nm�Ӌ�?k!��y��)�ע�M�C�B�b^[	�Us�KӒq�5���-�3��;m���%�˫�fk.h���	*�/%�JF^ZGR��]ͩr8_M3cI2�&�w�yp;	�v%p��.Ā�/Oo�i��w0���o�F��:��W~^m����_�6�2o��'K�j��!4)�~���H_v�V��W��}�w �:�C4L1�ّ�m��fu/c�?o�:�+�_��Q�T�t���4Yme��}m}\�b�U��\�g+��z���o�֎�������1xH���3�Z�u���{p�� �Q�=8doKc��M�C�?ݳSM����X}��ڒ~�'p;&��c���`n�)����W�fR�U�:���gR�a!$���4�9�T���G�r��Tu4�ڛ߹ tR
���;cjO������boE�d��*�d��Y[�}�$��S��<+�?�X�Obt��b�vh~E�MeN���5Y��e�����v�#�nlw�Dy0�י�n/��UV۷0�v�j\[�p�8���8.U��j�L�]�'�D k�澚��G���+�DČ
�����,#���JZ��S{;�_�9xʋ�3�z`ݒ���|����%VQ'����j��4T��^$8iۥ�fQ�7W�A������)S @�eZ{Y
���a��˄�g�O�O�5L�C3���������tJ�aT��NJs�=���F��H��oJ��N��>�0��P�(����w����7�|��x�(p��� ��#����QK���e��ςt;�r�K9�囋�EOOM��|:����fPB�$���=������@�����֫f>k����1�:D��i�sQʾc����������M��<:ŀv��DAk7�I�p�k}=⁎�A������\����F�Y�D���#�����%����!����F,EZ��{i��<����я��~�H;*zЮ(�mZ�zM��'s�}�3{���b��z2�̙��D�։������>��d��@C%�AΛ֊(W��էcή�N]/&�Ƒ9jB�Ǒi��0��Q-h��[���������+�o��]�kUzOc�z�xi�vL����k�NK�Z�~KpC�_>?"�u�5��u��gߩ;J�/mT���b�ҁ���ʗ&�]��Z�M���N����i�MUt�t?����Sc)Io��R����&91H+��4y�����|�&�1L�o���T$�U45��v�T*GԡLӎlӱ*۶�㰆=��{Y5<��9�N~[�?]����N��d��5�t�Z�3Q�Y�f��۪�7�W��[MWS���	��Ƣ_̎rp*��+ހ�7;���Cy'��zo؂$JN�P���c�_e%e�7U�%�zҏ=уd�5Â��`%�����	"�Ս�3��	��'�x)�b��+��K��r�|2�o�a��d���̍�ƴ����5(}`^n����@�p�#�����u.,��W>�XRx����ϧB0���C�Xy���?5.�X5�U�d��.��i�x�v88��mtY+�0��o�
F�f2*���{����d/u��<\s�^D6�-Н87�گ�b	D�1��U���u��R�gɆ�EY��ӱ(]�|=Q�\�&���W�l|$2�F3ò$B�_�~Mk�]� c˟��VtG
�?UF��s�	������^+;ܶ�	�@p4���?Mj�Vt��z���`3}ᔼ�6�M���F������/}w�0�s?��z3֍����rw�Ȁ:"���*�~&B$�F��?Nq5@��u�\�C�j�a�g�f[������aـe��L/#o�no+��/����ф�?s��)'oX���֟���:��<�LP�}�A�m6h5���z|���Zz�YE���R05?��?��+�7M��$�{�������u�-����e��?H�7Ou�b<ֺۉٚ��[�ZԌC3���y�|���sP�3�7T(�ؒTq�{���-��X ����M��E3������g��H�bR�K�+C�.�h�{�XT%i�a����[�e/d�>Tv�J��-
��lpv�%V�*��Z��3���$�13ڹ�}��})����ſQ�Eg�J/�Vj���8���J�+��p���8����5A�➻��S���X�����k�yV���B]�����1�!ПK�".�з���(тپ||kVw���@�!���v�M�$��{>��R��A��WN!�M��$ۖJϣ<����e�!֖j������v���ʏ�A?/�t�3��f���ٸ^���ȩ����HO�I����GW KU�䦰��.�������$����!M�K��hGc���U���\#��@nM\�qt�8�9�7x�K���Y��m�%h"�-3V�b7���-�������5�D]���B+��*5��"aa�N�D��/>��)��1U黨㥿�	m�Ţz�\��$I�G�M��=���uw&u�d�9e�+ܜ�y��kO�w��m!feSyШ`R*HKo1����:/�����}��8L��Ch|�����c�R��"�F	g�=z�̊�e��{W��ܐ�씒�:t��1�W0��]P��珱��fYȯ��l�ZC| ;�,Z1½>ɜD���*�I1�12��Pqo��8!T�>p��8��V��u���;�H�##�	K>�+�f�ÿ�2���qe`���b�WC�܆�5�׋����deA�!�cю����D�V]'_��%��.)J�����C��7�MB-�9{�F��M��h����C�����vz���ɔ���U��ٹ!�"��Ss�R�ta��]�������u�z��r`����[�W��Cs���_N�w�,�k��]M�-����y�U3�C�.yn�]����Po^�{-��d�m0�ݩ�k�鮕 ��Qu�%k�pǀx��)L�)�%�60�u�Me��o�^0�e1 햂�N�$������v�s�
�P3 �D1]�a��	�[3������O��I��Q5�M�)S��[,��R�x�U��H$HY~�p5��?�;B�k��ؒC�ζ���~_b��U��';>n<,��S;�_҅��,�#k#�0}WdiNu�C8��m%��)��韡T�(�h�H�~~Z[[�[ɍ�6�;����������2��Y�IKњ�F��m*�֎�<K��2vM��n��P��.�3�����39��S�	���&�;���H\o�&΅�uU�'w�"(s=��+��p��|Q{O;Q�x�-,4S��HA�n��Uxk��b��㉺�(5Mߊ���٘������դO�6��!<A3d�z��`��:����f��i8`E눞�����G_7�9b���r}	Mn���s8�z���wN��|*�\=�n{w�*�w�Lu<zD�"0\[(o)n��/?��`���K>���@$d?�����F�ʾ��Y��9�����>��m�$���LOb%��9ښ�9���h7z����~b�Qx�!����9y�����۩TrՄ+���L���IFSy�\�*�ԙ�)��sV�kh>ɚں���o�oY1�c���9ȴ�����+�!���z���.��߸$s�un��=ng&���[_�CϏ�#�mlP�\P���s�rf��sU+KL@x�?���s��
O��CZh3�;�e���É��]c��1�PFhw��_�����l~4��N��R��Gl����%w�C�,��v+�7�ac2푆#��^F7^��>ָ*�b�ug�j_:���I ��H��u4�$������e�����Z��U�Uq�l8��eܯ���������r	[�'���D��E���jE��}�G��?Y'�8��B��ǲV��E���J$�}�ỠK�Z�#o�HPM���m{3m'�W���"��i�����mj��iOI�o�OӋ�ⓐ����}�k�w�Jh���v�;���{C��bd$YyQ�w�q�Q2f�)����JD!�\sH���[�#p.�΅���¶g&����B�(�3�Q��v=���F^����?w���?G�Ed(2O�g�d�O�T���=2c/&��}p^�}�.ص�u��>���_�ª �	z���QRr�^/F�X���5^5��,�Y��57��r-�J\n=�H��p�xX�W�N��
��h-��]Wt��`�L�ah�����F۹�uH�o/������\]9!eǢ�^�0��*=�ܹ�����=�L��+
�k����������=���X`�t�=��Z�M��]���9�+��6'����-[p�`��!,���R��@�s3x(X�~��Z^��v�~���rkon��Æ�yK}�o���I�q-��҄4�gS<��8D�+�d�h�{�^�����z�7'v~�S��bIjtXf&#3 ��z�x�j,*�"�n2w��p�8��q����< �o���Zɤ���	 p�-��v窳���A�
�*��%�_�A���e�|�̜z����N��^��8~�'����iÂ3:m$��&�z��B|u 5NZ�7))7�z=V8�6>��j��^��& �9����IE��9�`vh.��:.@���{�ʗ���/'9f�!�[����6�*�ڋ}x�ޮ����ǧ�y6m w�11(E�
�輩��֒$���t2��BB>+_���gKsU�u�moޤ�� >�B�A
&^�nD@��6��UC�q��n���Zߐa!f��8�����=k�bV
��
[��HI�Ӳd`oM���!_Ժ������s�+�|�d�R�e˧��CC+
���n,�����ښn*ֶ�mֈ�B.�Z��T���#!k����PIFx�5���.���͑a��;I�YDpp�Ǹ�#K��_}j�8ۈ���#�K^�P�4vm�f&�<n�1�"��]�������W�CU���d�R�8�FF��X�G�ɬ��|���H�N�j|�ML�<A���!�Ϧ1���`�*g}�*��s�6��\�f�Jblx������	��K�.��-�=B8��X뷫A
w����-�8�g]���f�5b�{K����KG�'���K�>�i��1WSB�#o3�U*�� ���|s��u[n�=���Y?f�ɍ�����/��.���{�&�	od��}�^/���=u�vEZ�?�c�^Ȑ*HiF�ɪ��X�M
x ����)�]�dQe�gggs1�����<`Μ}��G��*)��1r��h>
(&t%Rd-k��<d��.��>l;�մƨ\e��?Z�Q�=�A��WǝܮL�(��k˟y�0_{�P���ٝu���ݞ,���nV���ol���?	��#�xk�t��w�g-�y3O����]x�<��;�r�q>���!y�4��Q�MЫ�P2��\���6�,�&� �:p�665-�HR
�Z����2s�p~��� �Ә2w��= "�zq�I	��3eEĲ����>L�cX{s���d<_"�s�Ll����#jx��.���F�u�"<�Hӗ4��Ȁ$v��T�8[Z
�""�����:]�o�(gϷ�}��z׸������t��yޥ��y�v��b�$֚=�p+��PW���Q)�ȇ ?_W'T]��d󏁳n<�v�	5���:_�>y;�^��ʛ��V��O���|vX�[4��[��Q�;�g$��	�9���;�e��w��ߢw�n�K�˻c�!�<�Gv�����g����l�,��سr��ʿ�%O�R�Zk�cq!��-8�U��E��|����I��x'��2�ϲ0R9|9�� ���e��}��v�/�������mǗ@~�q�l�%�<ٕF!៘ۜ��p�y8`u�+�3wib� A9i�K�L~	[}�(��ʆ�JD��wo��,P�Y�H@�����|i����2S�FS%鳫[�f� �j�5����`��he��ҥs�$*��F�����}.}��)���׳c��������[�yn��Ϸ
v�'0�*ole��?��8����<�J��?��9'�բ�-_�HF9�R`b�OEnw!����:�9�<���mz�S�%�����+(�U)�.-���9��A%|��(<,V��.�HG<���UX<�����iKYqW�n�8P@  �nTS!�A�k��I�l�C]�{4�U�EA$o�w���t��t�����L<��4c�Z�ϭ/��ľ��(�lL��@�����5�܎D��p���X]��6t�>|�������
rG��Z���������?l�<����w�"A���(w�gf�~�A{�D��nE=�hm�$I��o8V�v�S���������{�]#̝�Y#�9@.�2�̎EQ�d�V[��Юp�/���?����Q.?,�#����t�2�U���\��d9E)��#�v]vI�6��2�H0Q�f�}��Mi����݃-)�&il��q`k���516�SB��l����Q�t�h��Ĕ��/Ǌ��N���3�/ Gpw���LHi��l�{v^~��;��� �<�wD"��F��A���g���?���I�H)N�g(�� ���[̀�^~J���.D����䙀�ۗg�G.�9s�$��C��E�a\�4�q��M��E�hr}����[*�_����^�+�Q��
UǢ�7��!g�a�q���Je��5�>4v+����ũ�x|�r$�I���3M�]V~�d��,頙|�����I���?W�g�� ����F���!��Fa:�#'��*�&��S7ej�>�58����kN(�R۵.�>�o�3Y~s�_S'� �7�N�r����=�P���ej/�v��Vs	^�T����ya�q+��М����L��>A���اr�m0����^|'�T'���:���/�K������jJêk�4d�kLN����^QQ��WhP��b�_��o�ŸM�6&Ʈ�6w�C�2��[	5���{)o��t����)�����i���2��e�}�J����Y4H�&a�F��R�@��MQ��_Z��d������~�v���@�X����Z���@Z����~#Z�2��W�*<f̗��:-���
"+�Y���z����Ը��-��N�`3GԌ��U�뫙�Z��ȱ�8Q�w���~:���WM�#������B���u�ˎ��r��ŊQ�t�ԥEѥ!�i�&�)6���5l���XN��k�N���5��H�v��`��k�Σ�'�({D�c{�|*��'ުu�Z�u�n>�H��WO�I�R�ӛ`���x*���A�\u;!QɁ��K%������0���ScHyԓ�I�������������xiS�r�v�Y_�,�<]�7p��`����Ȝ�Q���'�L0�qnq^�sa})��M=���7RO��N�� ]��U�2/?��dKxȺ�WMXc�h5�~s˯����Ɔ�bA���v'qg��������k{���:��
�>����|�2�_NfWE|+����U��hs���\�	�A�L<O5�D�p:�w��i��y�0 �Q��l�*��*����	��֑O�fo��Ŝq�g~�c�3���sYۃ�j
��ż<�v��~��#Hh����f�y��� Я�d�"y��	"k�,[!�c��
��0��d�d�ROǽ�P�:����@\�(��a-��[�/�kF�ۋ�<eP�L=�ņ'Gёv����"�{ˡ:ⳤ4�q�c:&��^�Yp)�Ħ����>����ԥG���L�y�����:�Kw���l벃q*N��lYA�4�Á���),��v����#�Tɲ�=�x:a��Zf!Ft<�	��]1j�U��6���n������ma^�$*z��cuhxF`ܤ��������53���-�b.T
o��h��/�ߦ��4g����:{����*�x�<]m�>-�G{�L��#�O�����c�"�Z*�Gqp������%`��88�|�\j$�Q��$��܎$[>?(�\�1����D�K������^y�[�x8z>l�f�Ӯn�"��dt�7��n`Z��W�.r��ʻ�鯪C�~���R�&�ۄ�9��Ӓ��ә���[a���CUy#���Yw���(5���f�K� ����_t��$/����kw��H�CX�͆S�{9y��t�'_8�PH�@�q�%�^Z�a>*"�vm�z���;D�78lD���\d�*l���Q��f�S��'���~��������d5���&�|_>H�����9L��e��U>��=m�GA�v�f_�ryNyS�v:e�͓�aj��&��qgg1�� �)OX�K��h��Ru���O�������;����R��������(���[��<��_~C>���&��tH=�Vp��
#WK�ǌK0���z��P<p�DiTg�,�T�^f)�:�:��1J�^ڸ ���:*+�L����è�Ee<K�*I������e�mc����β��5a���1L�e��7#*)E~%�R煵���s�I{��D�\%��Nx�j@&�Tn�)����J7�ʂ����%�f&�?qg'r��+5}(O�hr������یl�f�:�����~>n3uF��x��pW�ƶZ��1ZRsTHg,V )n!7���j�O�'.�ƴX�_�p���w0��^XE'�T��rX4 Z&�<;�O��:
9��b+�gI��q7Wx����>ao� g �8-�a��@��m�։�u\D�b(��wg������>F"6�հ>�׭?zĒd	;���b��(�,F7.&u�;!���j�|��X��c�ϻo�H��~�\�w$����ޝ�"eDe��}�,9��g�{�N���G=q:tȑ5��|ڴ
�& 4cAZ�4��5�Z�����i�J����>��w*�$�n�a�]��T�y^���E�������;>���j�hC#x�6���m��RG�_�e�>у;�[�_���O��КF8 Un�4\^��%=���p��x�T J_oE?�~Zܾ�WB��uz"h�������R���	��q*�g�G��{}�ѫeu?rdD�D��;5���0�C��=�~�����)�i^`�(��Êd�6 uf��*'��d;N.HKj�Ʈqp�����{F�����{
a)]�.�P�7�~��gKV	]�gb�n�t�g����*�]ov��n�����P{L���5��~c�P��I���h��!�~�t�iP���E8dW�O��n�Ae�Jb�1%g�k���~�#�k�!����Q�=v��� /��wDXM��q����|��/E�CR�>^n�O
��cN���>{1M�]�^$5
���0�4#1�,N�܄���G��i��o1��9!��Du5<.�p	�{fz��$RL�#�Q�B�m��W&wi?]�#�]����&�2D�7QuoL�h?B-�+8����P�nw�>uȮYE,���5�,�����w���m��~@����ċ�բ�R!�ڷ�^�q�O�C���%m]LQ2s�E�|Nݰ�:�cSԻ3�[,������1:��^�u`QkpH[�ڂ�`����sD�2ͽ'����~	�Q�W��(��m
�hְ�މ�Z=C{� &1�aI�[{�H`f�����uSK�3��4*h��O�^1�����5��͹x��jp�Q�,�TUχr���� �Є��:zbW:�B�>��#��ˢ
@�=���]n^2D>�N�eu5sO��
~�:���.6a�4Ř�z��?4�|�R	[�!9����-Y^�B����Ei�.뼪	B�e�kQ�u���_�R��{ɴ"%�53��������ҤTg^�|3G������#�.��&
����| ��c�l�M��� �L牷 F�l�� ��}���i��d[A�\�kDۗ�Tki4EP�1��F�|��"�Uz��|����($|v#+j0%�z\�I%�E1�hoI��ɸHD�M��=�����Y�hpD(��[y� <1���Z|�����G)/�aʒ
0�w�� �6c�I˼���I3�)=�7ܯ 䝃�}[�����H�˻��gw��Ŏ(����<�q'Y��;a��ų�dY���Q�\3�������UO��!bvjxUȭQq��-����z�����/��Ԩ��e^�o#�R����L�}���5Z"���@����wOt!�	�p�%��ޡ-��f
�sU�NpQbQz��f�2��H��)��q�e1�6���'_a�Ӓi\r��D/�GG�������9��6A���9>� )d��0E��E��a�ڦ<E����������ߦ�':SO��A�̓����Pi�����[d5��da�����k_�lAlQCns����G�懠�y���J�T�PU\�o"AN��U͕(�W���NS��Ԏ���	a^=���D�}�+f�"w4�kD���n�{�Dd��&a��=���F0'��X���I��u�(�����WM� ��[�V=$�ۻ�.���h@Bd#�����ٱw�k*��X	k�w���g�yS���D�?5c)5�Q�i���=�����n��?V�Plz��$\�w�؝ܭ�B�5�kg8���E ��1V�cb)��[�S}����]%�y����� �5;e�����f�#l��y�B�q�k��6װ��r�*"(��n�VW��ܾvM�I��x^�4"?{~~(8EN�6��Y��2��z��,H�Zr�YN�����շ��F*GjEګ�n�����^���!��r��6A��^s���BY-��@���I{����w>�g�|oU��d�Dwsʈ�(�`Ū�v8����Ly��(�l⬻��H�&�B��Ks�H�bcFމ����Ɵɲ��S̒�BnFTE�p�n��ۥD��dZ"���������T&&�D�a_w�̀dݬy_o�%�O!e�GZ�4�cJH�  ^�!T��Lk�V���	{��mV�8(��?��G���8��Vgp�Wj�LnK�ي��w�-���C��>}��i�9w1�.���g|��,��9���,��<����{�ޕ��M��By]�ݟww�:��_n���
r��~aB�j=0w0��K��e�q@�_����X� y}�Qpۮ��C��m�6�_`e�+
�a�h`�I�^���֚��}�_�
�d�i(E�i���e��G��m}��B�֘�>wz"���i0v�kfWH�#���Q2�ߔ&P >(�AؗI����Y�_ W+;���vC��ܲ���J���a��@#~��,ە�Q�f'�?���~X���u����%0�!�y���Ƌ�9:�M�r:8v�{�5Z�d�b�qڴT�#x���A��W�WKL��btm��b[s{�(��tr8+~�����0��?���@�.��������������p&�{�v�Пv�L�;����X�t�Ȃ�㥼�@盱!�a��ge�-�!Y���Œ/S�z��~vo�:]�2��d�k!��0�@�oM}�ʯ��E�[0=ßj$��I��:+Q n@(As�4-Y����]���T�J��W��vD����feX|��v<UĂ+�Hk̶�tU��-��˹��K�yOdv�����j���Uϲ�i����Y�F�(�#��'=R|���)x��5�F,���j�X�ծT�׃ZR�z6���~z��iλC�*tX�E���g�t��Ei��0��m)�4�}5v�%��m�qs�3���ӄ�p�|�¬?�Wk��������T��b������)�>���`&���Y�N���X�N �4�����iE~����4�F_����24���uB��)W�;�i_��o���R��Ga0m�w
�Q�aч<1mڜ��3�{~}JM(�i���c��E���P�N�q8���Ɨ%�ȂKў'Hr�p4��=����ݿ}�Md�^CY���X���`���J����9�)���!�ȴ������W<stQ��V�I'IHQ<�a��g��ϻ�������>�B爻��tY_&����~;�N�PL��NJ�i�i��ഋ1�όA�Tr=���̄�9�;��L\�����O�{�gvW���U;W;��'f6���_x���t�ś;�_BоO�l�60���Vr������i<]s/B�I�lY<�O�<�l.��(5л�4���a���3�j�a�J�Scba����w��
A`�fjR_*<�W#3gpu�R<4����_&>lP��B>�	K�E(���I�j��$����@�7>�����ۏ�3A�Y�8���h-����в~Ij�#���`ھrF<��m�]�nƄ׳���:��̊-��2=�����5z��+�ئ^�;��~� 9��6�b]'���&��C���<��5�����;iSw�����1}����==֨�cOz�ݸL�Aa�{L���,a���x<��y�y���f���������`ȅ��+�Sa]���T�{f�ɮ�q���� lŃ��ήe:C�3Єvdh�J2χ  ��&��ˉ艆��["�^3�$ (���\@u�;R���И@�=`N�s>[k�����q�"�?���A��g���{j���Q�3����~�̽4?-�F�	��,܌�A�N��E>~�Cق9��2N��a��w�T���<c���1b���6V�aႨ��h�]A�D~�����������:�|!�(�0���w#���[۫)m�v�M��Ȫ��=���5�DD}��"��UB���0"M(���R��$�����ϫ*8zJ�"N'mEo@����`D�`{2+ �F��dJX]�Y�t7��`��}�{Y�µi ��C��ㅥ��fѡoW����}�
F�~�ĝ�u��g��v3���{߄��N�r�Rw)�֖�;zB�]�|��Wa��sCPl@�8�4�@��V�]I�#�Bf��k2�u��~��H�K�𕚬|����K��ӝB����&���cӖ�:�ఖ�nc̸8����"� ~���v����
i~�4���6l�3Z�b�a�˼��a��8٫��9�8�]�"���*lLf!�e���OT§�h�|7��Mc��I�* �Z
�s�(Jz���%�6=�sR_��s�̨�J"�#F����j'���-�_b�sh�F���]!U3 �1.� �!��x�mu�u�M^�&��PBA�6�Z�X��R���s_��ξָ�O���Hi#�{��9q�V�S"6o)~�b]f�	__'_uR_�����5QLB�4��=���;kĖ�P�p�쭅��&���h�h���ܦTV	�_L�e���5��E��rr�p���R�����8yӷ��ı<��V9�`͚��	|����T��E�k󿥃f�2V�����{D߳�T3W�f�FV�F&��e��ps4�Gn�Z�������0�]�5P�P9���B��P�P
�Ϭv}vH0���E�&�4E�Nʕ�\k����_1�ir<�h� \q[8)��P @�if�����WL�Gx��48)�*7��ԗ.���Q������av�y���e~��:;����N�_���}1��էfž>��!�;��§a����%��L��N1Lh�F��1>
�`��r��1)�]����x8`���l�F[���_̱�ԋ/��?P�kA##�-'/�����K�N�5�  Gz�nA�p"I !��h�<��cs����X��Q�BoQD���(�d���C¨�ոh-)��G���c�0r�b��q�ƶ�F,�C����&29=��U'��y<5F�+A�n���;24b������JT��B��i��H���R�����z�2���|��C� 9������XV(�f;]��������Š�>]����O�!�oE��ui�6ѥ�sZ�V��#�G=�P%&'<Q2�d�����b)*�@q��E ���//)=S�M�TG�$�S[�@<� {��co��皝����J�ߍ�Z\(�F(5�&�]�M���,X���~S�ܖ����k'���<e�H�a����_4����Tc���YҦ��4H0�y�l�(�E6	����E���J��Z��%����ͭ�ˏ��
5��ʸ���5���q,�yI����rk�(\�XC�C�4Vߕp�����R�R4�c0�C�&�w�m��#��/&�#�N$O�v셭N�Nb-�ι֍�����j̢H�[(�$e���P:H.�!S&�S�1�߭>�pq��G�d`lrF>�ᨫl����֥����Hm4E4N�ߊXC�,�ҁ"�iH$�q���-n���2x�]���$Yki��W�^v.��=`�}Ї]�~\�"�!�9鉣UA?����V�Qr����%��5�"�1��[��Qc�q�7�	�E�նSk�iI�8����5f;���G�ƾf6�\� ��Q��nK��3 	&:�0����;��BlK�aH)�����D��Ѡ�$�kR���s�h�,a{zn��m-�O9���έ�@���xi��$���D��		Ѹ�o��-dڏ���b)F�+k�5�gX��8���N�tq��R;	V֢�9F.ЧVya���S��5ٙ�����d�u,�:K�ڽ��0~Q}�����MrI��ߤĒz�ĝl 5q8p���OKbli��i�)��g6�e�G4���Z�i�c��F�E�L3W�����HЄRYSC5���On�`�#�E��*F4�8D����E:P[A��E���M�FA��d	��]�C�D�G���;l�	����`'�PV&9����	S�J.�r���+f9�Pq��c)���Ay�D��'^�����Xa�s>&4��BxE�q����g�DN)��%նdG�X���m���}�@���&ͪ����)s?�b���h�����O�ƍ�����ߝ��'�4�t#�I��	Ɩ�e�����Ź�_��{|ك�|�2�?cYdG_=�j�)Р z��)yk'q�(QuӅ���(Y��i�xbq�.΢B��7�R����Z���R��%3e�+6�h~�D��KaZQ�|�]��G�0N�W����Y� -�*>=N1�Q.ݞR�����b�x{�kG`8�L�.hA�Վ�d�2ы,���=��0>�ɘ^-<���l~�)<��AʗClu�J/�h���kO��/<���1�N83�#5_K���I.��kv|����Ы���8�ZNϪ2��K��Y;c�ƺ�mR
����%��7�N0�ѕV��!Ғ8�j0r�w�
��3��bI��Y�	�*ԍ��(�
3.����8��&���C^�V��L
tCLO-��POQ�kgvڪ�_�rX�'`5�OC"5Զ~IW����E��[)�/�Px85�,VL!��V��D�E��N����_q�f�F�7R���<$��n0�- �jߙ&2���{��LH	J�j��	�h�G�+��4^���?�`��j�,J5�����y�'���m%��|#��=��w�L��N���d>4!�<á���U'E�4i����!��-���+_�Є���'u�ʿ%��ִ�M�
��ʳ�@�#M�����<�&p��1*��ᑰ�~蹍ћ�E[���ʁq�5c��é;����ǃ��^��"�Df,s�P��O�Ab���j�)�Qs��VT>�	ȁV�����XyciH����JU	;�{V��{��s��>H���H��sV_TW	*����XA��.2Z�������w�B"�0������z��t5���(o��OHd � ����c�j�y^���r�f�jr׳�:�$*V�?�?Z��Bz���ϵ��������:'süW��G��w�x�����N�6|Lm|�ㅔ���A�_|���.<��0�]��s��h*7,#��XsDB��*�3�5͖	��t��]�٧
2��V��V I��?��2(έ�>		ndp������m����.���	��.�>8������)j��{����{@s<(�%ws�͐�=�;9\�<��h༻&JZ�&�T�rJLS����@�ʗ�^Wca��2�g���jrr��\�� �=�D�%��ti��E�s�(!+�e٠���2��y�;J1M�_ƁUYu�؇���%u�^���l���q_��h;�\�D��N���n�/s�ŸԻ��}�����-��B���Є�
!(�����N��y>�#y�r�b�2�D�NE��b����c��#e��]�G��$�f�e@\e��L#�|r���h�@�V~R�n��v/Ҋrb@ۭ�`fw,�UC�fu���uP:�gҁ"�e�n�ٟ�#�g��ֈ�eE�w�	f$�jJм|�Ȃ��) %J�_�~���we\��ˊ����0��P���;m�W�U1�L�ƾ�c�|�f��%��կL�L��^�AP͠hD��B+��_4��'��w��.j�ڼ�[c�?��s28����ؚ:�Ä�I���.���,0۷���p�	G3ttt:x]Dg�d�r{lI�Q1B���l��%*�>�V(�����+��H���S�.#��Q2�]�Z�]0˄��n刞�S����B%�I��yYt�Xt����td��o��; �5���
��;.�-2�lS)c�QY���Q S����jR0�PL�m9h�XCj�����=��R�9#.m����;$������K3p�g6^�Z�3c���
��/�|��7����
#(M)m�nq��`�5��K��@�l�_�F����D�H��F`?�~�t�"�/�� ���12�d�MG��(���i�@^eL��aC�s��3�]�)B���o��>�|�̞nϮ�����b��iΘk'�L�~]���͜�f�L�?63���{��@�%\�jr� ���p�V�a`:�c%Hi��5�ߡ��)�!1^S:��_�/�:��3I�������ͅK6͘����\�轚]�(`k�w�';�y8]	�]{�gW����+�f���;V?���00�E��A�ĂJ
dN�<���\���h u�{���]��B[b�f��x����0Ѩ}ע��];�M�k�N������������������:�7�Hd=W�{��[\S�m|��/2��h��n$��HYdWbK�t���	�2���ꁱ^����r����B��W$k���t�ߎ�$��y*���2^����r��[���~�;�)]�BI�!H�"�5?�������hߘH�-�8Yt�y���.�?$!W�G[!�޳=���3u]f�`�*c��|7�w
�6��e�=���T�uS�6vb6��>�
60��������ӨmI)��˧0F#��*��7뱋0c�X�c4i��BO.dJ�~�Ѻ�eZ�,$2_F���g�?����~`w���wuU��$���6>�.�(f�bp��
�A:����<�g�J2�-��M��ZnUgc�O���p�VW�6X�"y�C��}p3�P�>��㠥h���л���g�|�ܶ�LT�@OB_�7���1@fy���?�E����N���K�&�嚯�y��F��qX�P�8K��O���S�`	\ϴ��(�UT,��N�k��-a��c����Z�G����j��3��iK�)Ѽ�Q�~���m��ͭ��F���(�����zJ2�G"�"�r�%�Tm�Z���B�ɷz�ɨ�Dw=y�yޚf�3frn�%Xq<�Q.�&f1TR�CA��Y"��0h��(���r'ֺ���� fbQ��n���A��:�F��b����F�m�/�o���i$'F�9@'�O���#�`iA�������c����pqO����Q1(d�Û(%5��֣�`�7���9�����F�bha5��>Q�"��@�a֖�U�-O�F�)ĳ�k���'Y���O�&?���w�U��RZF��AxXY<WaU�wQs��/��Y���x�w��s���2h����-�����T���mc��/䅼��(w�*��A��!���#\}�wP�Gӕ�<"�'��8�H�Y��z9�iv�h��,y]����!Ę�c59-b3Ӎۖ�&Gt�F]4��/<�|
�VQ�yj�ղƴ�'sYm��;�'��w�c�U��琸����
?�x(��u��s���1|�8	Z5q�p�YIli+feF���8Yk �9_!��ƙ���a
�'@j���>�jl�#P��5��jL���)��fc~eRr�.W��6$��b�T���q����C��mw{��E�}�G���CL��~jBI<�\�_#�J��ܨ���a�2@I�Ws���}c6����Oz+3�ٱ1��~�Q[YHF�uLI��(���=O��7m}�I�]ƀY]��K�U�X��7�l��(�複��_b��9I�4kn�f]��R��1�Qn/�q�Dz��8��!����;ȯhB<���B�k�Ye.��{`>q�Ǒs9O$�с��F��Y�%�[5]x�8�������W�F�g	���l9�SG�QZ����#й�Fy4�IV�_��,����T;)���u��p�;�o*�I�1F�sȕȃ��a���$l���[�D�mL��uW�2h���B�k�I��]/���I辌�-�Ȇ��s-Q��S'-���I��0-m���a6AB�u�r�LF���Y�[�6�ת���z��AkK�kjĴ�oYR�ͿK.�uZC��&�������G�9Y�o�*�5��!����Q��x���Bw����Lj�jM�QI�z��\m+Μ>W�cA)�#�!_�麣s�*�,�;�ϗC�ʰ�G/gձ�b2��X����(8k���~#u8�	��(�L�0Egu�{?��]�]}�i|zɸ�rs���R8��:v�40�=Ju�x���7{�k�zg5��ߎ���)_�n�b�}K���o������զK2���ti�.=Y�#�tͳU�w �3}|T�1Rl��w�u��AŒ{r���d����F����\S�-s��UjV�ۓ���ɬu46�>:�����>c�{jT���U�]���j�����)í���.;�N̍�<Ӯ$���o�2��R:+�*b�ŘMߎC�XGm�Pzdb|ϓB.���Z4IG�"d�f��zىq����x���щ�R�j�C�*u'P�a����.�7G���">��c����_��	���&փ�O@�m�L����<5\Y�p��i�tO��� (��ڳږs�g��*}�a!��v���r"T����_AX0�oe�2�D�bAǰq�/���&���[%te8p���Y�As���?�k!]�}T
��Y�2�����(t����F��m����Wɨԕ��]F��mu�dR�u�V�a�G�PU%ΰ�!����
�BS@C� !)"��?���g#G/ݑS��.�br���0իe�圲gyN�of[ϣ@�d�Q�!�w��JZ_�[�@I[�o♪4�?b���[.YE���*x���%s��l8�
�8��[=�xZ��U�=EDD,����U��p�m�X�ۘ��j���:Ҋ��$ʨ6�.&Ab�}���._�N�${�w6��:���%Y4��L�����x�i%�va�U xA�/���`@�en��u��D��tь|��M����R|g<G�z�/��߾-xf,|�X�� ��'t���Y��F ���ݏø�8o��,��������	���e��V:uϖ�=���<��B��(�ޝ�=��W)u$�^���:$��b�UHQ���:�s�'�up?�����Gڡ�׃�dm����,�"������#�+�e ~�})�*�!y���?g��G}�s��Ñ),�)�Ѷ���|R:#-���	�5��yn�Ѻ�AM���UX{wjc���V?��2yn�Ϭo�Mthw�Lh��QYS�9�i�^4.�q�$��z4���i�Ŗ�����V����F���X�ߣ�h@G��7��5Ŭ%F�RՕ��6�Y�is��Ӧ�o]�;�}��u��9����͍��	1��bK�yg�C;WЩFA��>�Zw�=Zu��~�4[Y�ԣ\�c�`a�`����፶'|��K�53NȨ�Cr��^�7k�>�+�g�~��ve�t�7MJ��s��7jFQF<>Հ�PR��-�)jT���������/#�/�1�z��'|ءG+fhȒ&����}3�a0�^�����7������g�x�ÌK�e	̱=�tm���%�|��_Ϊ-qV��s��V;���OSG&������	�6l��qj¦�Ϝ~a�\���\�.��^ƈ䒌 M�;3S��O��K�M#1��q��G��~�c���Y/�Е9�*;��k�V��e���C,+��/W�9C��)���{&���ی�b����39/z��2�A���su�utQ�����@S��X#����N�����y:��/H@g�ƃra�_�8��_Э�t�F��d���f�稆��$R eT��K�:=�^��3�N��s����O��j�F���'�jJ�ENIM���YY%�#�Ǒ�R���kp�IFN��,�C�R���_��ۛ�U��� '�qeːM�n�~��Ӻ(�g\R�p�Ͽ���9�-س�88�y=�|�����ܫ��c�� }/��Ǖ �[�4��q�= >�����@�2~�*�iUu�yx�yD��4P�,ՋnJ%md�q�_�v���ʯ�I7��/��>�M�V0�+�1������f-J2��\���7�@`$e~��[�88�ʃ-��a�u�l<�&��>s�bk��=�����1z6�f��R{�(��o>M-�,-Y;+7�b)�A���0䎔�)$��+��\�,ꒄ�a���jKp��䕊9�����p9(_ȥ�c
�v�l�9S9�e�6/R*Mf��~��B\L��-hY@��P�b�+�X\��l({���eV��������y:�l���>��(7w�]N$`�9�Y���9.�#]ဖ���v_���6��U��_�/���-�C�"�ZWS%*P|�cN�9"�f�㵶�sF0\������b;��C������z6��$���^��_�8=���[[|�"$꒮���g�'|rۈ��xP� 9gs<P�涥ߒJ�}��
#�"�*�gU�#ꏑ��z��7"TFA>9bw���U�gt���4٩�ԅ$�AG��,�*/#:�����̾�ޏPt�L�u��z5��}���OR*8r>V�yFh�IRi�)�C'4��篐�H��t�x��2���F���&�hޯ�����YC�q��e[IX~��t
4���J��Y����Aq�Н2����p�����*��%��ώ���&m���-Z�]���]��*�l"_ �KS��������G�vJ�g7ݦ,�g��;GA�kQe�+/xV�"۵y���K��?�O�p�Pa(q���5ϓ���n�[\��~�X����<���
��*b��LdIm	�gd9�б9��ꏞT�_��eekjjL�V\zP�};�u�!�XC(����v1q��<I��ik��X^�qd����:w�1�d���Ĝ�y]_S���;��|�%H�/N�u&af�վ�C���B���UYZ"l���e���[�ڟ�tf)-Q��#��n&����G����ԼgѼC ����8���	����]YK>oX�Y���Ļ
!�Z��h%M� ���Zjj��%��޻�<R3z�l�gݪ��9���=�\���r՛hbڨ�0��:��ТܢL�t��Ίc{��1B��`��ib�"Lu��^,�����
�|�){쐵��F6�1!�<�j�I.�X�۾��Y��-�'��n��?��!����lJ`>��d���ƴy0*O8�2���<�&b�F�FS�i�b�#=�B��k�B9��c��ʿ���t���j�Ef_rU1�5��uZ&;,�k{PJK��ɫ$_�Yڇ�7�Z����6z���݃�|�@a~a�����DIRi��Z,$u�_4׋���Э�,�,a�����r�������zc6j���fBe���%Z�x�܊�O-��K!6��G�T��Sf��93��<%����Ih�j��Ex�����T��|�JLXE�����V]�޲��	���a�L� V��E���Rx�VC^I_j��&�Ֆ�ZU�1(ГE{��λ��J��V��ўMUisȢ��-��6��"�����&F+_��P���a=A�D��W�s�2�!�klX�d+S��L�Ec�ȿ���l'�zC4�lF5�f�{X1�%������X��=n�g�� ~�ׁʪ�k�.;�E�����Z��sVu2`s7�G��~t�B+&�`����/�l��~��;sYT�o��{H*wvk�o��:���i������ E��煎&x�6,���1����WA�/��V�����D4���A\E��t�r�#ؗ�`p�!����Ũ6Ag���$���+{��#s���F���޳@����>#���q����3HT�n�6��憔�>��qS�͈�;���;H~��Q%�hb��<~�7w]���b�dy�㖦���l�J��7g����s�E�FM(��H�(u��88�R���_G�>V��?z]@x�7��WZ�������+�u�g�)�X-<�.>m��F���-;��s?V:�!�l�OD�d�4�_hd>�0�n�\;q��dZ�[Pj ��|��/���bo9����
!�G*<r![*<��8q~�C[���'�^���3g����.�qN�G~>ЦQ�)G\;��S{t�AC$6=WuF4���)�b�{��@�i����_���O� �cfd�5���TSˑ�C�0�-�H-�����.b�/��a�ʺfԹ�X��F�?޻��`|����|`^6�%:^!0�v��	r�*��a�wL�<؉zv7��7�F�=)!�+�؟����ɝf�k}L�[_#���א��@���X��e(b�r'��m���;Y����B-g۔�Z�aӋ&����/�̜��Gj�EO@�(�m)�ߗ�I�F҉�I�c/����7�ki&�iDd9��6?�|#
���G�N��<�2����O��怫�u��s����J������]�${��''.��ahB�uE��!C�K�O����?��_�Y��Jk+���!e�	��q�蝒-�u�(��Q,kgZ%k�
֔�[�FLdK���ԎMkӼ[��Un�S
C{P�5D�鍊���j��̃ƛ��{e�� $���i"�n"�_c�]��r2rˤSC�}�t�)�V�[.�������M�_��n��B?e7>R6F$e���f#�2�`"�-'S�U�5!����k�+ڈOZ�4�|[W�	���e�m\��At������7��0�(��T�cI��5�*Qd�Bo���>�ܝ
��Fr�O/[��b�Y%�f����jw��+���թa�+�Ov��!^��j�P�
tٲig{��~0ؗ���_�4D-yr�d`�>���P�¼��*��T��t��;Y/zS�[�i�9����h�X��*�ww�H.�9-l,�<B�C8��N�+��k�^�Y%^�%^�|Lkv|A|����Ǘ����W{�G`�s�6�D-f���7�S|�{�K������K�����C��.v��#��Z�Ĺ����`:	��!붻o��9���1��A��lq���[ٵ����PE�`<rG�(E�^Ϥ0�7���AϳYn��L�b�@��)_-�KɊD�h�c�!K�c��:��Y��ns%�b�S��yM�9�#\�6�5z�2�>SGc/���7��ӝ�f��IK��#�oY{�O�X�s"Dp��|��(T���Zh��ՙ�9��E���;
��!�Gp[���95k��uj��:b~j�Oe{40�MF��;M�A��I��r8t�!u Jh~*�Y]�A����i��La�M����������Dۓ����ö��Uk�cf�X m�\�b��}f}jj4OG�(?������3R��PoD��c�W�Ω�O}?Y�_��3�꾊n�*���cY���K��9��)��#������-3�;�SbN��3J�:�u��U(�JW�}��ҌᙩSu�EHz�q�+ا���;���p�$/˰�&~��2��Q˵j`��n�{؜=n��*!�MW���
���\G�
�;T,S�*l)���4���h�NUه��)�Cqs�h뜔�O+�o�-4����15;4X��q�Ȧ�CN��p�,�K��)Q����/�����آ�#06?1���0h�-��y�F�n#�^Q�r��Tw�Obu==h;Θ:ͣ�"�>:�Z[:��1H%%]���W���<p�"�G�\n�@s��	�����' ��K������F��,����b�"��cȻ����*�f���R	~��b@aoP��������ܑSF�"4.�3|`׃�M�/�>>�ߊJc�����]w�@�怩AQ8�hJ�s'FP���z�3�^����<Wۗp�
RvX��IA��#���R�EY��dUcm�Ue��+i�d�H߅�@A�D9=IAο2F̜~;o�eU4V
�� �U����4��~7����2��R��=�ƕ�3z:}Ha���J����&c���J�Gtˏ�{̪��3���]^���B������b��{Ns4o+q��K����spF�5��ln�`c0��B��1���4��H�{��X��cX�Ĵ/ʶ�h�O���Jse(ܿs�$R��/'T��W)��G8�S���?*Լt<<�2=���;��;��լ4��p+���*�e���&7N����!�qs���Է3��B���K�����jŀ�#��+c���n�0#�ڢ���iX¶��׹���}1��q|�ϔ�/�$�!����U��4�Y2w��ٝ�� )6��������ӵ3�\hi 9�T���~��C��.�?�1$�)���[�?Z�UQ^��4U|.29����w�*P�I����!R�g�Iob���53\�������J�L�OCƘ�D��\$ z̗G���c������)��E�V�%�r\�z��_�xk
?q�ș�b�Ϯ/FO��}x��}4�O�eH���c����� #'|r���3��Z�3���Όs�k��'����?�򱱲
����1i{���a�aFJ�:R��@آ9�u�q�;è|F��7 .z)`�Ҝ�b:f��6^�@m}��}S�iV��O2�B
ٞgeH*ܚ�F�S���I�-d5�/�2���r���P�3�SuV�Ö,�w�Ї���P�b(*�uX��zr|ǝ]܊�k�h�q_>��<^�Nk�R�h�N؅f���G�M',Yj�V)����֐��g�����7����/��	�)
�1���~��;�����q��NB*���N-=�A���KfZ2�?��ț��;n��B���S�n�}0����#s󓇊P1�ZX����?��.���T�,y	������-Nvp�����8��Ia�� � �߲o����=Z�4F09��m1A39�o��ݔ"|�x/qg���)_��m9q:�����5������	���_	��]z��=
l6<H�!Q2����m��_�>
C�(���=�-�rR�y��8�ǖ]gkѯ7����{�h�Zq����<c�?N�20��*��e�G6���r3��@Z>;eQ���^�r��pu�7�g�dw�d�QÈ�?�Ǉ�Ae+��2��K>��`�
�Re--Qq�}���}��E�Ǟ<%���jjH�t��@�K��^�9��ꍜ	
R��GT�xV��_�W^�3��@�䍜�8��}��1�?���K���\%�&o�釱х����I��9M�գ�Qك���/W:yŚ҄���}9��Q��L�����}�$�'-7�и���1ںT'յ]�Ű�4�~[�{�Nb���c���d"���>�&?�Cn��bt\��V�;|�k_%y�2����*��!b+���)�/|��&լ 얟ńb�M[{�����7 ��$G��É���:oj�n����
�ͱQ5�E5�t�,�Y�l�%M������PXG$Bѱ��a�]Ζ�0��-�{���v�,"����s`�0Ly�R�N�7ׅd⸛��o��3s�bؖG�j�8�ߩ:#`���o���g�KQ�\_Q���D�ә����u�/2�t`n�a�����w��@����
\�`��RI8?t��U����q��,��-O�������J���L?��[������92s�!���;?�[���.�Iz�OA��5pv�L^J�N(G6k	�¶GK�9/x�K.��-����e�#�B�LX�xUYlT�����C����	'%
v,��r�$p�����m�'����Q�{�!e�(=Kd����R��'y8�-s�NvQVG4��r<��x��*3�x_�s�x>M+��]��v�����.r o9F{S>J��q�jv��o*����ö��������*<���5wl�Z.��2�jooN��B��H��}+ݼ��C�v��NC]oE��B��
���v��G̑f�
~����F�i�|����&DV��oG�v=z�}M�#��L�Ϊ��F<�o������\u���0~d���zJ�K?��e`���8��H��Oj�t�"Տ���)�EHK��vD����������R
��+��L���JE��P��)+S+���s�`�}�����k���������������&�1�̶?ӷ����a���i;q�G�M��p`-����Y[��Sf]`�J䝝˄�m���k��<Nn�4�����g���zUI˺�:yvӍ������1!��{���>?����Pݸ�#��rwe@��G"��p�{��
~�N�v�DNb2�nG�޳������(�_Y�c�.��⍪@}��:w�5��>O�0Z�ͅ	l�)�bl�����Fb�����C�?��1ˌ���+h��k�b_�ć�Sw�_# �8m3y>䳺6H���n5�F7��ػqϞ� C(O�7�$����CS6X>m^��^ϭ�~P������ީ �!]��#���kM^�����>�^�<�����r'A��m��/�z��q\2�W7K��q�O"�&��V)q�-��z?}y�湤m�������|�y�Cb��R!]�n���mݗ�eg��D'ӥI���Z֛��2�����bغQ:}	��ĦY��{(v�����XO^t�L�㜴��{T3�Q�>>��;zJ!�*(�O���o�ҍ�(��ed�e:���Z��[m�ӰUG���.���u��V�>5�ng	x%1#��PV�0��6���6�j��V��P�����x�8Fj��ֆ��{�B�^Sd�N�m��W;�M�ڎ�0�����m˼
�Pgم��6��&�8~��8���U��U�}k��HgW�6��q���/t$ڥ���H��F�$-u�L[��/�i����7������6�Y�|c�(9�#IW9����e�r�f���2��0ל�䖊�0�hV0��;�9�uZ�ȸ��p_�x� fhS�k�1r�.z���/���3�=������}
�eL9������l34@p-W���Ӛn|��L 'O5�12J�I� ��gk]�ʳ�ꚰ���^�s�<�Kn��B�<��|����P.�7k�����rg���W��x�|��N>�"�K'A �[@��{Λ{	=�:
�����baZRF��+�e��n����)��h������͍����x���b<-����E߂"�u�G�ۊ�vOsaV�d�^�ڋ��ltqD���Bf��nd��7ڡ��k�6�kz,���[�{Y��f/�]�04�ۇ�i~Gܬm��פ<��@�B&W㈜m㝍�V���%�3N��+W�,1�!~aѕ��m0�v|��s���:��[y*۵�gn]����n��^��1m:�A�_��`������/?�[pt���ðE0k�6;��g��^�w_`�{�D�Gn��m�NM�m���c>�W�C������HCv�X{�ܞ/v�Σ����f	$����s_��_x� 5��p�U��H~���2�+\�'�nD��T�R`l[����d�g�՚���rq�>�����2wh �24I�{�\l�d���x�#RB�R�ݶ7�8�����t��CH;˲�b�^�B�/�E��X;�Zr	8o�oK�GI��uc���OH?�8N���ָ��ƹ� mR�z����'"a픐�jq����,C�R�}ӃG�x1F�_�G�$��x���B���C=�z�us)Fs(F;',���& g�Xۂ�i�;�P�5z��.�{�{"���i�^|��#���m�R��;Oay��m^:J��x��;�7]�0)J����!ϛ��* ��/���j�CC�婢P��l��1�.�W|�� ��P[`���i�_�X�"��g`�:y%���77�^e���<I��-I�� >�����Q��{Rt�T��I6�ɖ#H�t��2F�.ߐ���5�Ęj��?yB>���ҍfbƚr��F�1�Y��;������4�6���fWh��m��j2�W9�28�{"M�Ct�t9Ȱ��p��"ņY$UZ:�oEC����)Ҩ��!t���(F~�"�}*X臉?��ĩ�?�4�Un,O��������X��Ip%k=���tS���_3���9�M#��E(�%)6�}���>�M������ޝїM�y6�l�n�T7֟T��_~�n>1޴3^����i����4xh^��韶 �3R^|,�K��6�K�{a�� �0�;|R�O��V��(����P٣�!ۏ��`=�M���-�<`S�G��3Z[)�����O�	N�JMÒ���;\���� �;G�?[?#g�Q��T3٥�=�����:����=����̇������U���Z���݋��I6>�V/z��T�����!�=���f8J�����l}Ho��i���M�v����a��5���E_n4?j��+�NTF�K��8/ޣ{}�=�ԋcBT�����y4�BA��1�S��ӑY�������P�+۝�ц[W�f�y\�
�ο�H���?��귻\a7W��5�l��It����+�t��bs��f�
 ��\(7��Ⱥ��ӑ����@מ�Vѩ���"C�����6�����Mv�\׈V��O��{-g�Ź{Z�p�ۈ�*����+����!�O<M)-�KtBQ�b���a����탉�u�u戋J<�8������IWd���v�?������4e���D2}������h$����_���+��T%-l�E,>�d=h0�X��e����V�*@�cV�S�V䤳G��v�Z��!���0�5�n�ϥ�<���ժy�L9�F�l^�؋lK��iU{�XǺy��~2�����:�����Q3-�l�Q��һ�����VfLsYԼ���4j���S����X�4��VK����Z��r�YmH��lna�Z1��������k� �-��۽��� ��Ñ�y��? ���{N�F�X����_i ���Y�4�/c]$�L��X���p��m��@�H��\9� A+G�:��!A�\�FFw���$���l���	����>����x!G�h�ԑC�&6ܕ_E*]�ę� ��#.�(4����q�?h���m�v��s����2�T�ĭ�������N��\���[��F�9���A�U¶�(n��cXV�0J=w���1�t����6���y�е����o��������0L۩�dʎ��䈋�sL��f�L��8~���?�8s��f2Q�
�Z�$�D�VY-�9��l(��*	ؒ�G�������#(�=b��ۥ0~�t�3���ڰ���">F�T�҂�1Q���|�H����^�L�C��MV'����IT�7�k����T>w��L΍�)����>G�����
��sY�R�%{[ ��7���#-�Sʂ�_jw����{	*�Rn�u�{�c��udN����9~�J�Y<�Vlo����dC�h�ůo�8*G#�p+�ً9�5N}�|��v8j�xVI��J�v�I�L�޶	#�Pe����dtrf�J!$rP���Z�!�T?�H8�(�$����A�o�\�5̫g�`Ȣ�� �q���FD��_���h���	r�ud9We�oXz�]��O6��{]�����s����[�?g�VvPa	7��Na��k�^�8��aM���
��rB�2���o&k�iy��6=+���Uo�������"�ɑ~ۘ��������q��-M��A�/H���YyH}�aK���S,?�h���{�C���>(0�62�q�����Q&��P �-$��i�ns�����u��r���%���,��i��PX��[�$J���c�Q����9��R�7?�	$�^�xu
qe�a����4�������O�B����b�o�W!p"=�=||m��؈0'�������SD�5E0�|G^�}��0R)�T���B4���ǭe���Oc��?��a� �_dOڱ��k�Vn5(8uS��r�:yG���d�����O��R�Uf+�Z魆?���"}��I b��p����^�\E�4���h�O2��N@�deI���qO֝~������w�_���������ᱛ9%[�|�4�[8�hEq���Y�ߘu��*�� �ݔ!�QJ�"�N�w�.?=�Z�u��P���gp;)D�����3�Xm|*���HJS���(h`��8�����E+�[�2��6L�1@3!����Y�#yȨ��v���N�XA�F��Z�q�^�r= ����ϳ�������	�K���3�&�w��k�=o�FDw	|�O=w!8{���\Ӈ��+�tN��y��?���x�E%��D���
�2R*=�����d�_6����H�doOe��ވe"z�7����8nh����
���!�L;�-*��An���j�/����mh�Y��Zm2�R�u���"LY�>��j���bv؇���!">I�o:��eI����Fד��k8ȣ>DKX"w�4��hx0�}��TD�(���]��>"G��^�U����������?��G
����
0���d7K빇�����2�bh�6���&��M�O3��I;���s���q_v�{����Ȉ�[��ʳ�$KjnC�>��k��[Mw�uj1xk�oߝ�c��3�s������ge{��I��9��B��;�w�ej�D�a�O��G@�A���5�t�Y��
���7�*J~�ڜ�����U/��������r�#�=��bR��v_�J�����D���=���QD�	)��SC ����j��]�!ﴭ.Z�v`�C�p�ef�[&K�>)e#Ff�f��W
�m-BUs8f�,SmS2x���c���ܽi����������ۛ�j9ɮ/r�U8ma�^p?�4��6��v	�ܪ>³'��[ �1e_Q���z�UBs{J��à����tZ?�W�=�W2]��$��c���ȳ>��������d���� �I#b?=ά�����c^�!�����N����d �^�bP��y�B�/Ƀ�0����g<5)�����Z-Z2���CW�@ ��Ҥ�9U�_u��F?(�E�ݬ/��?.&;�gSݤ�섉a���y��r�� ǽ�q��`GF��V�}R���N�,h�rT�!��)�W�;�!2w[�Yǣn+8Z��Օ���$s%lZ�/�����]�}��?�g�1k�Nh�Iҿf7@�����C@��ޔZ�|>���� 
����k�����s��d��)S���A�!��a�� �ǀ!���HUӴVN�<���q�샩H�%}�w�_��'3�BխV���C�g�ɣd�� � 胴�����r	*�9�G�}��6�W����q}�M6�rfMDs{]s�Xvpu�B�g��B�4<�l�/գg��l�!p�/d���_�����>ȑC�9:�� �/pc:՞�E����06?�=�*�}��j�6�a��t �U���|׶|����}w��?Ԕ,������q��1�A�W�����	�e8ݔ7���G�r�R*�����2���GW{[�dT���b���4i���u:��G�`�3%�k��)���BIo���ś�b���V(�_CF2����$a����'%J/JG�Lk�4
���'%�|wB��tT�kpA��oчɉ��[���-Y�"��Q�&x0�%|���5�Kѧf5`����Y�[�����X��˙�!/�`������
��Tx!fP�T�A�È�
�2����sͼ�Oð8����w��r���%�vS]��I ��-� ե3��e�;�#Ý���UT\]�-�����5�Ɲ Ip�������!�;��qw�I~�ι�����z���*��j�,�R� �-�c�$���uUd��j:c�����1ƗC�%��~��f�w�����q�_�s������5e\~�;�GF+��t�I��D��M�y5j����8^
��=ۍ�~"���r���R8
KO��;���;�~m�}~�*������Y��R	�%��V۔Ϸ�I�\���,�@�KB�j��ދ-�ٖJ|�g���R�X\��'��M��P��?���cQm�&N���o/�WKv,=��H��S)�MI�l���ʹ�٘��۱�͉ϥ݄W �b�����w&+�r�"Xe �����_C���V}�v�m����jȂޛ�a_〖�._���r��'��}'�զ���d@4qf�wB��G�՞^���p '�c����y���n�l��P���g���{��Y��F�����3rJ�%�0�E��]ؑ>��1m���o�NhE�[���ɣ�V_�`=H�?�B�y�߂ؑĂ�t}f����@��_+o�UE�����A|� �5��-��"N��f��,In��#�����(�a�Z�	~z�Е��69cS����^^ׂ�ȋ���wنY3Q3��M�Vmy�ǲ	������?=/OJ��������f�c�tө���P�K4rP�ׯk�m�I�����'���01^�CC�Ud?��kV�bĪ{%f,�w;�:>vs�Z:HkF���2�����2	^�q�Q;�l�� ����y�[!���c�"�������4�S���N�h;KB�W�"�0}*��qH�6�����1�B��p�RK��q�+�PS��<��ɝ+��^)��4mBj����
֜����1����@�U��&܋35]�o��*@�����z�<e�=P�_��A��<܎!�M��VN�Z����>#U�5��l�/R��o?��i�j�h���τ9x>YQ{-R��Ѡ�H{�Hj��h~4��$�Qj5�m��������L����|õ�4W\��x�S�ql�#�H4��߃��s�T�km$�[no��z�:!�wg���5�n���9�:7��˩��֤h���D�\��_cA��œI��3�8�$l�&�!%��E�X��q�ekN�I�D���h�qѵ}#L�����-h D ��xHk��{�ÖD�ę��R������֙�F[��WIw��ݭS�;��x�*3�����㖢c��I��^ȕ�H��b�'��Qx�[��n��-���Z�}U�E'c���6L�k�i큥rA�%�E�i����/��PR[|[n6X����ʕ��ؼ_�b6�{�^%����5.L`麽!���q�Vf΢�Ax<��hq�{7V��s#�Lp8�v���`hRe�}�3� �l'k
B�F֪&'M���]	JYx�K�v�z���-��0:XLPӭ��F�"�Dw�B/a����%LY����4��9�3��������Lሉ�R��.꼌������
�#u��b:$+�ڌ�7k=ok�	fv����,⻰,�L�l¤�=X(���W��A�2�p��ڢ�$�յ��?I�����f7�O/������Zѵ\���	m~_�֝�����!�p��w0ٮ�[/ܣ��T�Bﲸ����߃��Q�W���7��̀�K/���bE�>��V+d��q��?�	�"��*�u%�_�'�������-&������|wl|���*a������@,�����え{��˕HT[�_�E#����%CW{���gg&C�.�l�k��։���8�¹�"��D�$\�������ރzߺZ�XC�F���IN��3�8?Յ���ޟ�D�O���[��I_uڏ��m�e�KZo����i�;�kd��k+�L���$Z+Qo��r��v�IO�wP�[b��י�s5������Л��<*����'�H0
`c)�lzw��v�����<�=�b��]���q�I��s�i�U}?�}L�NF���=�UAA��Ц��ݎ�cCU'R%`���1�ع���3�+v/�l�𒫺zr-��|8��+b���K_���ɒwSl�:l�_^j	NW-�2x��2�m�����p�Gm���a��'�1�|5��v����9 �I�;����I�<�����￺ً�I8s�f��y������̝�X�;�1zo�������n���Nt,]4y �茳D��M�(�r�Ơ��;�O՟�ߧ��hu�Y_F4�C���Y��3�|� K,���%6z�βъ������-�X�6��<�e=E��X�h�f��W���I�����$�wk�&##�U�X��~瀏�������v<n3��Y�l�ۄ��<_چa�t��]'���-%y�B�:�&�2���itz�q��3��b ��C�c�{w�R��3��ąJo��i��Lũ5���2I\_<��IU����0/�$���dx�P�w%���l?#E���\�܄AQl�G�4��+�Wx��c+Q�މ�uw���E�z���]�%��Fq�O�ݹ�X�qv�z$��&$L�&��	���� ���=�����Tþ�3����-E\���Ȇ�u�;%,�L�L�U�y����ĉ�	饻n��{������cJȠ�7a�f<{��-c��&)��h"�g�>o|��
�� ��S��sc���D[���J��N��8Q^�k=А�`6׫[c8���+�<z��[9_�|�d��ߢ����AgDĈ�����*0L|gxNiU9�%��	V�<�l=9���V�m�ê%���m�F�x��������5�+�t��E܄����<,����оv�yz�U��ڰ��p��q�w�I0W�E�2���+j$�RC�`�/��i�t��n�������mRJ�O�j!&f{����BJ�g8D�v�O���dm�G>�f���.���5���g$��|\��˂�B|1��IʁA_,�B��@mO�.��������`ҫA\a!���>$"�L��l�~HY1�m�_��ɿ�BG%_�<�j��V������g�-�tMXx5e����A[�������;|�Ľ��!�@ٞ��V�ut+�z�����@o�(I�m�W�ID������qp�+r�v!�J�SX������5����GDDt�m�n�����@������Vs`˩�w��g���	"�u�,F�C8F��N˲�\CM�DK&0i��e2La�L��F�m,FJ�ŏ?}���P��B^�;�װw4�|��}܅E}�e1�.�Ľ��%$Ն3ZfS��=FB/|*F�qdw�,p-E���V�Q������"�i|��r��qm�ކ�g7������hv�Z4�u��jK�.���$j�'�@)h����A�JD��s��CL�.�����R5osf��]Ps����iBt���#��Xa�l�I��������~� uN�O'�oX-`g}���On��Q[0��
UsG>O-�m�E;xEU=8���>�5�64�(Xyh��7r�?8�[�7Ŀn�G��%��&��T�����Z�_ ��]�D���>c1�Y�*E�� �xg��Ħ�I�t3{`�Ǝ4��+]	�a@*��JV������a�G��b����_=��(��O�\ɩ��c+�h��E2�,�����ɀI��"�߸������b�kws����R�_ˡK��x�}�`yxt<y��nA�]B��ތ��4I�;WH�|=�f�v��������}7�?�����$�ng>��g����	�;qE� �A5�#f�GC���"+D_��[|C%C\nι>֊�>��= �	����8[���w�dK����9�l.<'f*����b��~=ӫ:B<_�{�!����q��H�����6_uKC�"�X6E%�W�j;����j!P�w0[��f�(��>�~���^�I�G_L_�8�<r68�(�����DW8El��_�}4�RX�~F�i\%@����sf3lM\�}�x:f�r����5=�/�_�U�P�Ii���5��#H�#O~;�<43��'Li��%��o��?�znM/�/��D��:8�G#�C� �V,Pv�P�d�EE���L��U�Jս��H�N�SFL���J 0��{�w�%���u%��,I9d�)�ˆ)�b���6�� ��+�!���U����n���o�5�qf�ڲ2���Pc`�KuBbe�F�lM1�������F�1�:���Bp��z����i��V$���P�_���с����s�¤�k��G1+�2Ɓ��2rTF�׷�9�B�]�s��]�<�%/��#�Nb�Ž�H�ӂ����;"���aPx�ag��B��V����y��&/ &��y���x�>��q�T�I��%M:��d7A=��8�#(zn�;L� �����
\�Q��P-H��ڗ�,����n�c�i������52=����'��� ��i�L�9�b�@�0��7����d����2*���QOG�.g(a��%�tقB�b�c�����O	-�Mv���H�v�
�vl{~o�P@.���g��l�2�i]񭠏!�*�M�@|jl��O���p�Ns��֦�\��n����!:[ǟ�H�	$��B��磉n��f�gX�[���:���M��|����^���x0;iJ�b�\�PX[m֍����t��z��d���[ػWI8���/zxZ��O/��E������p�,(RAA]-����8��M[< ���<��\�8�t�=�{����W)G��p;j2�OL?� ��+���Xjzw��^hRM��h}��`����ǘ.����`���B������g�D钼��/��=�:њT�1;}��HH��(^�+s-�%�	Z��E2���ՏV���Zu��J�Q��� s�X\v�*��F�`���C�Ud���|W+[ь�`.�� ����#|�8;�jev'�.�꼥�����)5L�T��RՠkWӞ��oW�*�x��j:*ca��ڲ���
i��ɡ�1�]5�t�:�\pO(�n{� ��J�j��:�~�d,Y�8ͬ�	A=��F���Zl���N���w���L�b��dC@���Q�{5h,��օ��D�W"�Qp���G|�a'�n(ߟ
x��SSu�R�ݽ�P�5%����p&�&Bhf�(�/���J)�A���.���~[d��(K,$�?M���z�Av�t
�Wt��n�b�����64pGW�g>�z
�𼊸܈x�?����B>����r�̊$�f� q{���"�E��#�$�鯟5��m�+q6{b��m!��׭�4ģ�V�_��#�_d
A��@M=S�tY�=��%)���0���+m�ӭMȇ��u�I~�򺿉*�r�`��Æ��R噾yxK��'���\%S޾�1p̰B��A�F#ﶕaQQ֓j=���>6�6HݰI�Pj����	�υRS���w����ɮ�&o�+�㎥���:oF�-�;�kz�.��m�׆m��>��'���Xm���6c���E��飏?Y�f�z���ʦ�Pb�NN���H)}q\�NqQ=��Z�C�B��t�|�ܭ�p��&L5�w*�h�`��TԿ&����}Xcho��?���hg+�U�'{�'o�1b+�������h�X�I������� �Y���K�(�dp��,���i���<�4�@.(�	F͵5j�64,��l�s��(�b� ��*�ڲ)���:�&A�>���ф$v�e|�5!H<|	��S��]=�y%�M�d�9y_�ֱ�{nuxs�b�-ͅ�BA�n�'��#S	>bԯ��s��*� �1�^���SG���!�G�/D����/UO�M�-)�aHA�`�^]�
�% �ֵ _��Y)��(Z�Q"D�b��S�����Y<hg�����'�6��3�/xz����/gԮJ?�-W��?��KI�z:�YG���5z�*���}zXp ��l�>�h�i��o5�Vҫ�����DG�ƿ�3�5u��`�� �E.�R=	�X��.O���qy��!*<F�Rf 7OprWR|+����K�e�h-�A�|�@"����`��۴0�63�ɋ���r�v����N�~&Y�/�ml��}�&�GC���(R�7;i�Gzv��*�4���S-�j&��]k�6u���c*4�n^n��[N�](X�J`ȡȣ<��'@gHݤ�J���-5�懨G*7`q��eSdg���~�ǟ����m���2_���؇"��{�BA�m�C����� 4��js�C˘|�}¼3�92K�+lDV�W�4M��t7怄�@���Q��O�D!�K��a���N����6:U�+�r.g�ʥ��dE�I�,Qϙ�yJm.�磌�L�uR (P�,G�i�FL�G3C[�g�6'@�������v�s�>�!/��'�{�I��H�VpS��A䬖�����BISP�@��/g`MR��،��|o.���J��b�N�`�l�B���Z�\��L��p���?��:KJ��䵈h
� UA���F|5��b����A�V�dDe��F�&p�`���y/����I�����y	16]�YI���z� /���^ܦ�����bۥ�4��5M�!�U�Q�6ɧ]o��)4��[Q���H����|`b�3(�.ͱ����-P,j�:��3Gh&�^�Q�z��3ܖ��/��+X�A��(9p�E�a��˪@��y����le�6�:>/w��-�x0zC997noQb�'��=��]��Ws��A��֢wY~��67�,sĸ��Fm.l"2z��L��p��҉��FL tEʽ��}��+�IP��Ym0g��Q�<�	q���ⶶ2���	�c�<������{���ٹ���U�Jՙf��p77��.v5���9Ҵ�F_��B�������#�oMQ�S�ىM���\}e�
;_wh�7��HL ���d��8T�;O�U�pLv/.(B~i���\>t�1�Ki�"�7�EDז�G�9j�a6��̦�_�]tFIx��C5�7Ϥ���a(.&��Gܸ���(��F�v{ۺ����"ӹ��n���	mD�˄�2���4�K�]�z�q#cѲ�-[A��,c�8��ά[�	x�I�<�u�qIjGS���e����`c������f+`
����˼��r�9}ry��ZD����`��uZ���p޶��1�l@���Jh��W69o����pB�{l�{�fk�r�����7~��\O�G���X�� �Dnp�;�:�\[ؗ$�ѱ�	a2�+��S�=%����⦫��+��2wTQ����9|��,��]j�������b	��������^����桁	��65Ã�zE���ѫM�?jy'��M���k�_�:U�f��yKv���Y.�\�ǡbd�6ԧ,�R���Fd�c�&��¢�qI�
����:�����"{}����0�L��F8��Mg�7����Vs����X)����S����#&��f��
���a��%���6!����������Y��NV�:5ֳ�a'O�Z%e���Bഴ��<���$��յi��"��d)��wW�~"q{�ҟ�<$Q6����U�֩���9t��ȯ-�$�d��`�ɺ+���<k���ԑz�g8�R�w@]/g�#�Rň,M!�B�/��8��n�w�<����P��(Aą�C��Or<�o~����
���׎��5��QF�8*o���x�~FCjt�3b ��֖�+�����g����퍏�˹�J���ƍ0�Ë�Oτkh_�����,#Wy�&���ߠf��R�;�����H��s}A�n;r�% �x�HR檪���E~{��(q� C�/W�3�����G(~���MМy�
�e�P���Ms��j��l �~r0wҷ��M{J��j�6��vv�Kc𲗅2]?�:�d(�\_��]��t�݂1��_c�*�V#�m4c���{.=��Ay�ZW�[�/?�g��v�ল��Zh�s5����J������������B�Q�� <�]%v�g���mY��/e8��͈�\k���u&�s&����?�?�l��q��~�ު�-�=!� 0�S�K���s BI�]��:�p�̖^1����7f3hzr}�ghc�+���S�Ϻ>2�8��e�������^:N3u�1:z7�*u_���4ۥ`ƞ&�XDi��#ߝ�e��'�x]w	\_�t���_��B|�@O�B����{�ȅ���z��Z�ր�9�5=� ���Y�Z�OҿN�wR���3�Y�Ђr�Ǚ�w�_�Hl�kvj�5��^�Y9Ɛ	�pY��/}�|����"B�7�m�'qiK�*���	[v�xOȞ,*C����|���.%UC�V~��$��E���3��~!��!��c��,��G�Fb��������њ�l{�y�z������CY7��!�I4!ɺ��� )�^S��at:ip�0���������#��NpUj�]������޼iB؜b�[#��v���I�b����������e}�w�,�?���������I'98.J��y����rkK�K����6�Dz��:it���+���x�_:t�z%B'��������d݁��ʵ�Z���iC�vM���e���s������ �� �Lڒ�Z��_�,�#|�4�i�ǚ�g�r1���:z�:�g�M̪�����($0�d~Q}A�3��9�5�%�.�� $�qx�hr�v���Ψ���RQ~��׉������MK���7�!��_!�_x�0#������K���F���0��� L�^7_���ݑ��}Q��u7�XY�3Y�8�_X�b��Zx���/<��p�:��׹o�<Pa��Y�7i���X�w��iS�Q� �cu	㡾\�(�G���O�K�� ������ۈ>5:�k�ݡ�=1�m|���3:]�R	�p~�z��y�X��C�g|~ȥ4�$*�km{a~��za�:���<��辑���ʖ�I?bm��h�I�/`K�[��F*�R��GŮaj�`A���t�z�Ŵ��)+�h������ks���{�N{�B8���U��u�wOF� _�e�I�J�Yd��7�ޔ�����m� ��5��Q�T-����]9VZ;����)� J�"c�,C��jT`�t�;�t�b$��@_snT(��C'r]����d�񆢵��Z�fqX-��-WK�,L$��^���I�����9�O��N�xckP]�Id�ãÔ��-}�A)�/���m���˘=�?�y{�^���;L}�U;���p�*�^�T60��|���4t/�5.T�*��鮿�	�>�h<縹��aF��{p���4eq�p̗۫&�"����,�f�8��Ŀ�:��"�f�`�Sz�6�B;�(, �K�m�'����JV���7a� {�-ڋm�k-�I�&���[.zv��\T����\��T�M��Gr������� K~J&}e�"�Z8�%v�q`2�h��:,�\&Q��&8^��w;fs��*6�~�S�l_��Ku�O|q�Q~����r���)�h�k��nE�ށޞ�@2/ΡG���F����u�8���6R���a;�ђ���z���Hլ��1�\�[S��ծ�1矮��p��ߞ�=+W{���,�+O5��؎,�{����� J��xd�Iu�w�>�5]�4$����S���sKJ��]�m�q��p^縉���Z�\�W�E��9H1�]�{<�I$�&��;Z�]�0X�{��;��V��a��$�8@Ax}���\Ӗ�ěW��������)�������;���$�A�"���\� �TkG� � "f�����Wq��2��HVpQB��T�n2�n��oob��G�I�!a^��S�"��6����"�`ɬ��ß�T��&D[3y�~��w3�x�p����аcr��z������ѧ���2Yi?,oLWn�l&�5�{!!�i������ց�I�>ͳU2�
�eti��d!�
$*��֡~��̀�n�������B��;6s�����4~���T݂iCw�Ϝ�[=�#�1��1/$�^�v��5x4�&�+%(;[�e�vC��CB���7���p�3RǍ�����4	8�6�����R<;K����Z��І��]Kz"�1��)�&�In��h�B0X�|nZ�q ���;p9�$b�ǚ�ձ��~�7����]
�m����w�p&�#�WV(S_����U`�N���',(ZH��N�yc�8 ������}���,�ed�_��u�#�
�����{�H�#Ҳj�eix];�ꬍ�{�Í~M�u=ҹ�rlѡ��[�Pu�>ן?�4 �i���>�i�����kkdRÜ�����s�n8�c:����c�.sv�ge�-	��<p�y{`�oyk#O�L�F8.�K�"�t�g�,Ðq���[����`�nܐ���7�I�Z� ��Ȥ�xk}fʃ��
R��+�:\���AI�JZHB�u|t�^���#~:Ώ�x�v�J��'p2;�lq��M���R}?�Y8�y�Cu'Jr::�TFKЌ{\{2J�"kF����N��H�T�P����;A����u^]0��~5
˓��c5�͎���o�㿁�Y{�ǆ��{�f��ʈ���%i��D"���I�I�6��
)=�>�pRt\�tyݿ�3R&�=�f��N��A�ˬt�^��6'Z^�2��72�dt���PO�Q���,�R�M��������XCk/���2S�ܹ)�:	f��@��9�c���Bu�������B^���cp%~XD��HsOȢȊ�E�md�L�0 �袋�L���K��ā�ٗ��s5���(�K�J�s6�QP��&x�7��"�-.��K@"���)g�C%��inE}"*}�������9���Y�}V���s� �!�L2�z-��/��䓩�-7$�窝���{�Pt��(��˗?3�l�>7�<uWE�<�ά�"���"���[Өc&ɣ��Ch!vai�{�ZQlE`�]��g�/��q�W� 2�SX��
T����F3g�'ȥ��]y;��⑪\a�aI�7(��@� ��5r���(d�G�G:b?6��~u$G�qVj�Cո���~�j�M���˿N|�&�_5Q̿t �*3s�ՠ���aH`婷�Mg�IHM7-�8�c��QKŀZ)xH�lҢ,A�8X�s�w=�fL�S���*+-�9�Pv<
U	���P��h��艠O�������7ޓ9��� oi.�EL�,K��.O L� �5"VW�|��cK�Nm@A�.��˲�-p�ȓ��	��3���w�+��(��.�d�A�Sf�-+ \���D"�Hy�S~o�;������2��׊,a=��������f����^�	���f��EG��?�qK˕ �3��ќB�!��u��%��@]�Lƃ�,�x�4��<��2���6�� =Z78b.9�/^o��>ѡ=(��zG�}�*�Ii.�܀I�m�+��b���.����ۺG�������kmؔ��o*Vv<�����.$הK��;�֏�%�q�������[д���3�]�|�+��d�4�7ח�ܽC_�T���+J��o�(����K��ɩ�q�K�~D\i��� �M%��8BD"��
�r�1S�z�I��k�k�Pi�!C7����ЛR�X)��`U�:��{Y�U�"�?�&�`@uF@��N�g�m���zU�a��a޺�Ę������\��M+㐬��D��0��Fk*��8�oe�9�A���`D	�̽?�|���pč��M=Q�ө<R]�q�cbT2&�|xZ2&:�K%�3��c"�~�[[��>D���hT�k&�AW�qŹ5�Xqg� ;v/� S}t�����D��Φ3)y�|�avL�C~�T��G��@gx";q�#v6�>�/�n����hi͑�}^0�J
��,��n�t벨%p��yx����Q4�}}.�֜�-�>�"�芲*�eOa;��>�Q���'���(�d�
H�@.>/����g̑���j�j|R��q#ٲϓ��<Vu����p�؁gu����_����4}��6�� �P�i�NӃ �BL�������St�꼂d�K��A���Gz�f����F�!�J�Uޟ���RI����[J��Ӝ�����Q�W�o�[Z�d�J p�3H��H�f[U�ڶ�[����E����+���Z�0�O���Tt��>]��+I� ����pS{z�����Y�R-Ԗ=�|I�&��,��3�}����jF*P��9�L�z��JH��-��/R}���p�V��+���J$���D�x��t���>��p��9��&�Y�Mv�����d��+��^�hC{�J��$�[�%ΦjK8���q��y��=� �Nč팁�h��Z��UD2y�.۝�|
E�{��K���{��o.���{OM��_�dBQtH�c��,	����C/%HoC����vS���;_��:���u��k�ϕ�����g��w����?J��n+
�{��+�[����Y��*]��dY��v�!{ޞ&w|�7���a��Pj�����d붒$\���m4��#?�Y���7 �p�_֟���P,��;y*ߘ13������M@�2"�N���@LC��G�	�	�M���C�F@�W��kZ�t�e����_e~;��\5)��"��.�j;*�l'�B=�u��w��3��~t�y�#F S	��U��
��;<
�_�`��F�������
�n2�O���jfh���w 9�|�8����}�)ѷx��؍9�q��������F{��[�W/I����vz�.���m��y_}1J�[�)�;l��@�x�jc�ȆoX1���i\�ČΖ�n����X��3�gp���95�2��{�~�<��_��7����a�Z��B��L�A���"_�Q"�Oc�����?�Z�P{zG�Q��������O5�L�&lzh�"QL�t����N�m��� g�D	J�CϵV,�I][4(��'�a�6�eu�Q�`sѱ�<E=񻷞/�㾡W
b�eN��/�ت�҂�e��]s��p9O~�����&+js�J�E�?x �+���-*�]��Q:r=f%�#����}����b?u�,�扳�?�h�S�[i�(����?Id	�)z�f����`zB��oy,��J2��^�ލ�7��1��nn��-�7X�����4�^�WVI���8�+��s�<��=x�~/��)x7��M�>�{g"5�3����!~�<:r�����X�����?��C�Z��1���H�,=�]������r�f�*-{��x�FF�ĕz"���$�V�Gڰ:��j�J���4��x��Y|�S%���ښ,��$m2�{�j�
=��ݴ���b��D�b�nJJ���`Up�,����[��UN�R��z�3�J;_���Ed�q�A�]*·E3\:B�pQ�艟eپ[l@�a��s�;���E�Q��3k��;��1Y������B���RS�{4td ����*I�Dt��Ƚ� 6�EGm�2&5/�m�1�Iٖ��9fU�=��= �Qm�ލ���ȇh6AD�l��nz����Y�o�*?�zW�"rX��iY�^x�F��93��,��3��S8#%CC��d�8�����e�Uo|ŮBY�)後�+��Yd<��Q�.�����G"�!ù!ZA�ֹ<�d�Q���w�	�Ó4��E|�UG�~in�@i`��v5��eh5��і�{��1q2�0����_�䲰���1��Z��)&Z�ѱ� Q3�g�b����9�^���=�]�[�Fk4�]Y��d�UT'�Hl| ]����$��53�������E�2�`"n� >*��,�+��4��_�e=�2j�K,�T0߮}xm5㟁�;-����P6G8��١b�ws�m��WvL�ֽ��R!�5����n�6@^�f�Wۢ�?��9��L(��֫u�Մ 3:���k��8ܸ�/��i��,SS�}�"��L�F%�?���۵�g���ڽʙ)]W0��zLWMCXu�;1U�$��=�	"1����T5�P�zٽZ�Zn�	XD����9���!k��# �::�W��wrglY�f:���a+�+��✛y2��YBb�L�'4�0h��K���D�y:gc�_;_R
tDd}5����5P@��_��:����~�ᥴ6!��vZ�Ty����׍�����%�f}fc&?������ΰ�� 4�H�9�/P�s�Ͽx�>�e�E����2��6OO�֪�>e�$qՄ�u)�n������~>�_^ʯ��2�A�}���NL���@2�B���j`C��,�I�V@��Zl���m:��-����wƚ&T�H�#�H;�����j�E;w�^�s�3G�վ+�'�2Ő�.���-��5��6Θ�U�n���#4벭
{��S��t�k'��o��{�;j��]~V����$^b����Ӑ2� z�W�+%�C#�_;�p}~��Z,�{O8`��º�x��<-O�<NYS����:Ԩ,ѣ1��>�s;� }����D=Kʹg{�-t>>��"����S����W����i�@G��u	��w������;�m��t;Mm�X������ RrY�6_�(L6p7�f��]9w�$=m����LUxS�g>�J���V�AK�w���֯���=l�M���;��D^�%%�3�
�	Om#ALAI�������>�ԖU4.���N��!���c`ʏ�Y����B���<��n�|�A��i[8���1a�����D����.�&�C'�*%�����sN����cڱ��~��N�Bޣ5
a�O�M���0Tl��&���q�����i>]���>.�>�]�u�֙��ӥhm]2{���[}}�n�x���+�$�C�+��"��-Sow���i��\�(��F���b�~^B�,q��fn��0 ҩ��,
8����!T�%d?���S�f�HN=3�X'jc��t��\AB����ȵZ�+��\�}M!��՟0�V�Z��A6��\^�����	��̾�k�N��!+~7/A����%�$\�'1�����<|Q�ٙ�em�{P�����0�z���.�+��+�Kj;s�[��<ɢ��]U����8B^A�NZ�VP��#eV��(�����=V�	R�ami��a��ԯ�7+(�fH��;���M��C�:��� �E�<�%�|�O��j�2[w����ˊ���Zm<^�(ݣf�rߚ	���r����o){"��^�F�rl����A���1qTpeY�;ޥg��)D����Q�>p�3��ז�jL��*�N��aMN�5ǋ{@5}�/Je��e��M��1zi0�Sn�2�h�Cа�O.A�<�+9&��L��𡮊�>��,��aP���0��'��L<�2���`��r��3U[��S�m��:\l�W�J�ē���>S��C�gM�,e���pX��2���w�|�|r����J� 3Q�μ��,g�h`
+;X.��u�H��k�e�/0;$�J�m ,��@Dx~��j�q��@	/w0	ʭ��ѫ7ҙ��ԕ4�@�Maݝ;�?xF�bh��*�����$&�*B,{	����gD�.潲���2��F.��n7]�R����Q���+�K]�_�05z:��>bb��f� #?��{���ܗ�U,g��g;'�zU#�e(\��#�g�Ć��r՗az���ٛF�$(m*�R��d�4�b�����2��t/"P�#Ky�Jr�m�{��%ݜ�+�n��t��߼�W��l���8e�4������05�^|�8p>%k��G��0��/������E�?躇9��з�.[K�@����ٶٻ)3 �4פ�OX�<%����M�lD���8�c��@����"�����~`]�sQ[f�����Y�,�R�n��
��!rfV�7���o			��g�<���<��Qe����\ٹ�'���H�� }�>7�4Ɇaϻ��K�A�"���՘��<> ��L6��	T��ii\��kޭ�Q�M��{����Ɠ��u�F�,\q�F_䃵 D_�ء���ޖ���p�7����L�3��|�Y�ʜ���nO�-v#�(��I�([����7��)pTL�|����kKv
x0@� �K1�m_����pg�ǥ똿OH��9���<�}��B�m������	Ζ>the�U�n(���t�ٕ��D4�.ι��e����.D�����,2831u�:��,�h0���火��:�3�x�љ��Ϩ3��ml���_��5�dg�0�f#�U���<�#s���#���K������D��Ã,���K�����z�8�`k4	������������	���A�������s׽�Z��x������},-Kbԯ��(4v��Pk�uy�g3�bygu�܃���a��〢_�ki�C�l�{�9��anu=e�Y,��W/e����h��3��7���{�D�	Dڈ�)-}��ʝ�x&�s�~�C��Y3�eY-+�dc�r}�U.oPkT�-x�v�M%î���s�>�%��f�4�	G3�'k��1f�Nm_���ϩG�ҖC�/���W17v�B�k-8���Z�AC�4i�a��n�����Ԍ��e4���慘6�9~���@$a��导:>S�Q��y���6Ȇb́UB��;.�<�o�@c�{��%.���<@��0Pg�_��ʈ�����,����"��o��\-U�ݭ���O��SM+�
w�~�OF!9R�3��+]�vy���a����'j�{�g�O�#c��{�v}'�����O�)�;��c�ki�^΢�tW�1��rf�z�
���wm5�����?h��ꥌFdPz\�9�뺤k����踑�">��0!Ae8noa��u�R��3�==����(�X��@��Ĳ��6����]`�*�[��y>�x�#�pն�;6�ݗ����P7����T N��KO?�~e���Ff`+F����Agm���/��мշ\G�%ɎU����BB����$�5ڑ����z��b��t��߱�Цm�)�X�YO�kS.�g��T\3�m�+��d_oT;�T��:��Q����P�*�Mwc����jk�M!z]3���P6lȦ��	Sg�vYZ>|z�mzQ�*�o��j�U�RY�>����%ãYsX}��[�\̢,�`��!���d�
���a���(�������̟���S�ج!H�Ī�ņ��&�ޒ-D;&뇿��wn�����s������*j�鐫�x�JήB|�%Ym��d��/�U�wٞ�y�T�ޚ��\��e�&C I#�ɘ]�?EL��{���f�x����<����o��p����>q��͈�u=����vSl�V�{�*��E��!�{#
���RJ-G�~��0��e(A{���y����79N��|�Nek���g��υ���T|����Mn���d{�X7�V���Y�?qގb^�M����P@<��ohܾ�ʃ�HI�+��W������HM1��e����xk�ہ�}|����0�}��h���7��(�'3�Z:��̸Ö�@�w�"��"�Q�s��wq�g��\'�
K�� ql�����}�>ʇL�l�F���RK�w���[8V;6��!��.�AP5O�����,>6�,���w��[�HW�M�8l� x�v�b��e�Eal��L�����D��V�:��؉y [�)Ge�q�i붯���ũ�f->Rm��-���~��p�9�o����6:<�8��q��������!������x�־ھͽV��W��ohOS�GE�"5�:ZW2��*���O@C�|�f�-��r����j�aOz��Vµ����P�/���N$*�ghhlʸxi�x�BK�!!����v
/��ܣ�li�y��XrK��5�r
)��u��k4'1�m�߳y��A�6�"^�'��GR��cl���.:��67���}�W�\�v��y(�f�Ӥ�v)�S3�WR��j+�66�| F1��mL���j��.��j�5��m#���f`�.�������l�\+��B�O���%�jfzk���o@un��P�@u�X�c��տ�E������Ջ^殂��6�N��o!"�ﭫF�ޞVu���D�JPL��]�뙪�p����%�Z�^���E�GL�x���<��.'��g����z1�5��&�Y 	{/cG{s���S���:����d�y�3��?���+^�Tچ�K��Ն������ET���2 ���s�! {�7��Ls�D��Lp*2(�o�f���,��9���e#�>�>���r��'k Vf�Fp��m�f7w��E5��]�Q�G��/��ꀿ����^�����o��-��\��h����.�C�gCK�ń���
��Н����R�T9�!(!����t"�⼆�D*���==�`�3�
��٣Xg��9	i!��O5Q/��!��^,����zoRͪhPS���7WT���_N�ΰW�s�0�%?�����!Kf�@�uT[�Kz	1���ڷe�lJl"�4sT;Ҏ�O�OC)$ih5~C�ގ��8�ŪR�(_5s/�>�3!3�ܨ��Q��`�k�����y�d�=�h΋��k�:4٦�SG��QYNK�oݾOX�˯��¡�d^�R��j��Z�5}�E�å��]$Tyy�A>�KI�Ųs~&ʩW�R�Z��5���+UG���Bo[����ӡ8.=�*Ix���G_��sf��}Smb?0gpe���t=�B�B�w$Vq���"��:o:�P�[�F�t���5��l-�pR�ͽ�K'Z�.�N�%�|�,͎	 ���Q��xq|^>ˢ,'���c6�9��\n�?��O�#^�x�$�Kn���J0���xd�kS c��O��z��\��O�=�5�e�L�7zj�S=J�8@����'`>E����fP{�9��G�M��b��_�X���Y1dD	A`J�PŻ�Ż�����z�j��F�_@d�C��E��l���� J �yy�7~�ٟ���~�P��}1,��v���ǁT���a /lG���ܛ�:���ol~7De΅!�){Rg\������(�$�<� >
f&�Zi���:�
)L����\��Sr=@{]^xrxC�2\"���t�~k��_��1(�3Cg��n~]�%ĝ>A�rb���<�d7��U\)5��!�n�,Gd$���Kʗ-1n���\z��lA�ha��@S���x\n���q��u��V���D���_����t�0!=f�A��E8R��e"��"�-N���oV*By۝��T��Mɉ*�s��7��r	@wZ��4N�R�Yv���{!ܤkZ�B��}�2�2k��'{�
���f�����[��~s�e��\�7K-I��]7')��v�����@Oܪϣ��u|}s��O%O���>��M�G�9�)e��7xV`�n�a�2�L��/�k��#N�V�PR��77��l��K�i� ��+������\	�N�YF�]�_��sV�I�	1N1�{�
��*������SK?s%��__G
u(W"q&,r�mey1E,�(k�2���%Ul�n��J������[���~4;���;�?ub�|p/r��=q��.�����Wf������i�K����h�*_+�@����N1�TT{ED��oN~�|���+��-F�?�hr�wr�eD�p���pC�_���Kr�@/��@��m4Ԡb���>�0���<klf�$Đ1�wʷ˩P��n���{~�iy�ة$V\N�jyH��LW�F�� QCScfE�k!B�6����gZGq]�-Y�0��Yg��/���k|�3V��?ͩ��W1�:;� O��ɭ ��>=��j�{��`F*�#=�b:� )uY4D����~3X���'@Y�q�4[���<T��'%���ckxD(��L�O�O����ƌ�A�)�Z2r�?���?����7ӷ$m��T�����.�����'9e$9i�u��c�*���dc�_#��&��@f�����Y�ߜ�h=�ԛڧ_1\Z˅���������(��|}�U����,�QG1p/O�0��jj�-)@<�x+�࿈�*��$�f�`���?J���H�P����Qw��okε4�:�QE���n��K=�5o��s�W�uD57[<��
��7'�v=�
 ��)�P�^g�����C&·��px9-f��WU��%C�$�*�M&�R��_�i�s{����(��>���	��� |׳��E,Q��������4v��i�ڭ��/��o�ym�������� Y��y���(���e7��f[� ��!�υ��[���^� #�	9�-�@2��3���ls<g�v�{Tl.�E(,�
�q�"�i��.��nz��ӏ�V➜�d�'�l�ҕz� ���2��?,��{�}/7��"]n[���\h���p��dQ�e�R"JYy�SR�1py�
�48>���KF���-̎E��y��~�?qG���O�D����M'�7Ves:��wZ�s:�"��9�q
Z%���\�_.�aV�s7�;E��9��8��4��]�l��zd��)��2��^Y��\3u	�+�DV��G���E�O��;}���Sq(�~F��}���s_i��'~z�����$V'�P~�2�rGu����4f dR��A=�0C�Q��)����Źz�j���w�I��W���E��j؜���Q�[����61QX�2i�-a�B� H��q~J%�e;����j�	kmr"���U��I�����!MZ~��V��ObVe���Hy�۪P�%�-�"q���A�US�+E]�U�6����I�a�HnE�=��9�E_�7rD���y��Ä�Vq����l�<p�n��	B^L?Ybn�7h�/���9���H��4~Mtx"�w��$�,<Wp)���M��&�*er�L��㋟��z��Vo�#l��2dSR��=pQ�
�{�H(��aq�� ewnyT�/&0UU��� �\�R�)}�*ϣ�䡗���S�lo{��5��%�Q��j��H�B��c����5�+�Eo����2����zFJ�rB���F�㷚ʩ"�Z�vY�\BJ�I+�TD=�T�c59-7�y�4U�8N�U'���ΐ�p�0�WR����Q[\��Ԏ���[�+E�%�Sd������}�bL�ˤ�9��VP 2�D���ȻϪ+�Ǫ9��PTS>��09��9��1��ɧ�6�ml#��ec�������ZK�մ�xT��Cϩd�P�Z�=���Nzgu���{4o9r�r}��?�!�H}괧J����M����/��;���(ߛ:$�_�ָQ4׽kj�"�LPV����'��"�n]�HO�����&��ѼB}P��ٷv������h�yW������h������2�Pȟz�.kœ��&7����X��-�c��Y��V�����
VL�Xl+���nk���Ұ=�a���޴�Q;xz�c��%s�&�o��R!q���8��E.ܝ��w��� ;ձ��/U�{��%:���`*^�Yr��<r�6��i��B	C/�>
 9�#s4pd��7?^���9﷤�i�B7Aێ��<��N9~n�I3&���jD��rb���j��<��JK�X��D�G��nD"�aL��i��}׋���x�����w�/>>eWjܒ�	NH�Npk�7�S��ϻ�l���d�6p���C�;o�>O�ZGGwx_T
��m%Ԟ}Tx.�����4�5���Pd2�Ȣg���$��v\M'MHG�3�ma��1F/i�D{D8x�3�̚�%�A΁�M��?�6���HV��`�uqH��j��UM��ɥ�1�����S�0ͣ��	!Q��P�{�%��C���$�Un��i_�heP�5��+� ��$��l�H�ݝ3L�<��� ��/�5������{�66��eI���*T{'�!�pR��T�*��P��Е�+$�_�$�H��:ԑ�����2�xE����З`v{�U��!�7Z�����;�>5��C�I��^�:N/1xmI+?�N��gË�e#(���[p�S�����D2�lH��x�Q̍�FBk��HWU>�����ݝX�&}���W�8��|�m�CQs_�Q�*�U�4�����Pʖ��cd>$�~:Z����l,1�J
�=�HZ�u|�u͹��ru���j;" V�x��.$hvPř&ĉ@�Iڐ� hÍ�]�XeODGI�4`2���4x�A+߰�g�.tI�����<A���AF1Y(7ܙ;L�(�ѣ��"u=��i�
K��K0?��;��9SɃT��p ��ۓ
0�.�I���BnN¤�����aX�j-x���Ʋ^?K�J��U�7.~Zo[���?  �ʞ -P�F�PْY(��%�-��v����O��^��u�g�za� �45�/>x,W�
�����7`j�{P������3��z��*Y
-a,m�@>�p+^�K?�ӵ4��z�Xܔ=���g	(�.��Hi+<��*����s�꿥������T�v � �ؾ�:�{��e"V�� �;$̾�L-���S�ԁ�	����J�,��� >q�]��� ���;ȸe���f^�x����3�PF��'B�.��������r���m�=�aIܴ�޻'�{�xj=����24�y�t؟a';�u��Vk<�9�v�t�[LZI,����cؖ��T7��&m.mӗ�v:�����C�m�H�Z?��sS����us$��Ը���.��1n@0t�W�s�hN)�MEx�n��H�(kBqBx�;dK�òބ�w|A�L��0���r��{�>.a���G G�1���f��=˲���;��H>pq�-d:���5����{$��
�O�h�+{ʘ�i�R���]�C�U���ZX[��%}�	�=h��� �k�o���c�$�6s��D�B�/z�-��r=g��~W���y��``�Rl���=�G�|a���|]T��|�hO-�>���>A�
���Cx�|����9�&x$�Y]R<n�(l��ۍ�0(*����W����9�й��6���)�%�6�͹�I�����#r:+��uK�O]Q[d����C��+�_��Wn���h{߯���d����좑�ntq��M��1_o��xsx}Y���)i�t��]��bl�{e�{�a�m�~�SE�;!�}�����Js�_�M �(7�T��4����u(�Ў�e(a��K7m���t��q���mx_����A6T��3t�}��քL�<_���8��Iq,�>��l��2BSy6�(�@'qH|�c��=-�q_mE���L��~%��%��v'^��\��.���A�7i�@gT:'S����l��U��'�Q_R�Sˠ� (�,�yJ�<�;I���>7�%�X�b�ݫ�#m��y`�<�O���0���a\#���~|�51�O�ywhw���5MxJ��?.)8ɰ�U�yf��䳒����L�tU�i(�U��6��3�h�EsL���5ۢK�ƒ��5�,��8
k�!⨕T_O�5�=��=Y+���]Y_On�օp)-S?���������z�����X�����ZȠ�إ�:�D�z��֎�#*�zBn�xB�a#2V}�?\�!Utcۂk�Y(���si8��E�����>�Y}�@LBYE���89�q&��@�g��C����0�_�c
��"q`!<���l���O+s2D����ȢJ��ua���0#K��#zT+�1������v������6Й�!�lw��~_.6Mӂ��6`h,E6.- W���c��"4J�M|��E G[L�<)�/��<�D��+�f��͠'(�V��(��X5f�]�<ԏٗ�;��QZAG�jз�0�á:D�ɦ�	���PX���0gZ���,:�h��|[��lAT�V�ՉĢ'H�(�A�P���n/�'*�Hq]�Ä���F�W��ԍ��+P�������"n��K�����-��o�.��"О:�4gA���-z�n�����i�qJ��c�8���}o�O�%�oF�۳&�VG��ɀ*2���ѷg��n�ZC�	&tl��&���aaV󰚞��0�$,]�	6��q��g��7.I����u���	M�����M{ϼ�ѯ�J�@}�:�"�1�T}���d�=�O��cD���j�	}x�"�o�O��Ci8y�b`����&��#��U��Vs��nךDL�ul吇\N�7?�ώ�!�u}C�}����B���F��_L%gm���Sy�jˊr��A �``Br#?�Hy�+�M��5��BC-�I'�D-ajSk��o���7����fs���mͦ汊��\c�8�c��{%��Q��gzj)�C��|���X4ǟ4CŌ���jy��.�Mo{��&�!�i�m/��5���Z�lG�t�b�so��'޶�c�� ͘_]��r����eW�~-|b�+A;T]�O�_�Ǿu(�<���E�����Ɂ-�� F�D9����c�,��`T��!c������]�I}b��{#B����C	�$��P�v� ���4V�(�ס�ˤS
`��H�7[���=��i0��J����i��Fn{�f�L�mp�T�d���j�eDFb)�1�����ɕe�a:�g�]��KSU�s�����h������(������[~ �0�T�M���<0?��oۉ��XdQ�Y6�f�`�*������"|ߋ���ē���2��c��Mx�adY���qN�5U�u(�3G���)��#ʹ"cꓴ?v���ޭXT	�-�	��K��1>�I�zirn�eD�^���OU=1��;�{��
s(��V���hT>C_($t�%��؊�ǿhKS�<�ߝq_Uf�/�� ��ۦ����$N�7�G"i�^\6p*0��։t�������/��{�½����?����,�����nX����ߜ=|�����"8cz5B���A���O�W��ՓG=>T�V��V����պF�y��m��g��Q#Ʋ1��3F�ݝ�T��~�~�^��OU#�|�H���eU����ӻؼ*2E:6�};�gΒ�<�rdG��E��o�x�nZ*��BG�cZ��+������_{gץ%pV�ݘ"m� �$𐥪��{_Qv�d��r�>����zM�c�jR�m������I�ը|�w�Z��ʉ��"��~���G7�@Ɍ�q���o?/����J�o���	g��B��o�q@N+XN�(�}Z���0�<��ȸ��R�z��O)���]f
�L�nl���)���$�$ͣy����A��R����֍��C�G�K���}d�UU��L�c���&}��M�!�����A{�;�������?�jS�s\Q��;p�������Ml�,f��q�b �Ý>�
ęZ]M��{�]�����1���OO`e>�<GP�\k#�X��f�ܛ�p,+_I�9�R+��5�ɼo�[��%6z�heޒW97|���lZ�M, �)0�(����5i.���ph,-�%P嚞��*7:*���;o�"�
-�W��������XBK��Ձ0T�0�$i���53?�ƴ��Ϧ������o�n9|wt*��o��ҼjO�����s�S�msng�+����3�Dܚ�p�#�O�����2�ӝ���C�/J�U'?�5���>��_��S�U����j�c�/&����2"tҶ������<j�t$�)�)1��?��凉��'�P�a���?N�Z��ݓ��� g)�L/�� ��h���kZG���w?���#K�݆�1���C���2-���:�
�U�XA���ֹ\��?y#fҜ�7����s��=+��yY�e���Fh�`��Rᝀ������~C�~2y(ʘ���!܀ZGl}���k9����n�Nt;!h:Y}*� �F�c�>�ڃ`��8\��+��&l���%��Iltxڔc������27�,vc{����yP&��6�a��++�ƞy����J��2�G��E���7�Ή��P���r�Tia�7�RT<���9v��_��	�l��,Ia�#*���з:��4��N*���G�ZR0�Hr"�)�U�:��ܤ��H���g�Ԡz"�t����ؙ�?�E쭻��l�H�$J�n��7��7�z�9��*��Y��p�R�x�^���fn�*W��#�R�7\�[sq���<WH�5ۍ �.�+�N�`Nb�)�e\
GYz�cU*�s���Y<]˧uk{fB���*��������������r�N ��4�y�oA0|�DFǉI�]���b���Y۰/������D��Ѷ�V5���Oʄ���pvCsg_2~����ܬ޶U<+�+�':�U�F������%G`���mp�v�R�p���l��U�Zr�w��ͣi{�����m�y���u�b�����ho7P��3�S�\p7�+��k	E�~2�	*���ea�:uKӋ��5����k?�<�"���ﮞKe���Q�>;	���*�91���<di5R}�dQ;����j�9x�E(��~���}�/z�L���)�a�I�3��	�U��H�aq�Z`"�-�L����|�U�&�y�yC2��Pz:�<{[T��`�};�^�HNI�X�������I�׎�����3럊�"m�0M����OuV���/@��)ܙ��!�Ģȋc�Ǵ��5>	��:������{C��k��M�g��s����};�E�eI޾e�U�;3����Zo�[�erQt�`�����jz�RF��bGS�r���&
��)r���_��ϒ����#����T���|���^}༄z4��=f��[i�(�/q�{�k��(����O}>�.8Xt�W��I�G�=4�d�]��U�m��^\�?���qnjx��W�.F���'�F~���ӧ���c+�����s�ξ�%�zn"Io\%��AS�e��jav]�3��Y_�
�Z:�(]�-�w閦�r��j�q\���PB�N�(3��"}&�~gV��y�Hc~�o<�>��ō
 C}m���^R��pԶ5��gǭ�����5��l��oU�'�i�x��Izx��o�y���f����卻PS0ˡL$u*҈�ts��K]Ml�Fq�;nĒG�9��#�O�^����)߸�(��v��[������X^]�'V�T�y����ʹ� ��H�L@r �ڲ/�J�X���[��2�i�I�	X'Q3)��vFqKJ9јoc���gZ�cM������B�@?��%Ω���^xD�7�Ѩ��׮��븟��e�v��� Mq��$	�&3�	��{6v>şO���:��-�*ǰ2��:=/���&a��n������}ş��/�1>Q�`jf7�7 2y������e0E��1��Q���ǰ�vh�7�ESg�����8��E�;'�X`��H��c� �`ϖ�M��9�*�G�1kŵ��O�W_��bBO$�v��u}��c�{�$���zM�9�HO�)��Q2.�ɨU�k2�� j����\vy��!��F��TA���d�/�l|}w�biRX�h��ܲ��6�;s���RO�v�o
6Į�(X�kIk��ԣ��@�̉X!��y�x,�)�Ƿr��#�t��7o�09��]���`7��Ŷ���$
0�=P������{�?[�S����Ob���{���fqt��[R����s.���F\�S+��wUV��(<̞��i'9S[���1��
E����c�����f0���D䮏�9ǵ�����ݜ}�I��ak
᳭�8�W�M@��������o��z��;����㟡��,;
���<I���ߪ���}[�� :qaw��l�S���_Ll�b��n �2͙�s��(z?(��La�C?A
]Y*IY���&W�I�C'>m�5����$x�TʞQ�z$Urx�26���/.L��'�:�������L�lA�1U����{L'S��A!���J(��*U��ܖ���� 5}�LF�y��?���#��?4�2Z�S�Р~��	ý~.�GR�[=�p[Q�%	!=��v+��_�wKT��T�b�ԧ8�e�7������T�,��
T�/����{S6���+��j^[���҅f��5yS//n��+���T���3r)�5$�7�+������?5;v������h
E�_�2��NbnIj��0oTb`=���X� �1�d�~Ԯq��,�#��V,�.U��A��&H��Gt��S������>DG�c�q��?��|S0U��Tv���f���u��Pc|��ru����tX|e����N?�K�q�0���{�bM������,��e2�+�ӌIS
é��f����n�&�p�]ژ��g��9�����~P�WY�?��a�*����R��r8���}�n�� .��{o�/~�����­��6�����#�6 ?���
~��XG$B"���Ǜ?�@�������}w��ǕB�9*��Q4ac���.+����=\ע����t��e|E��2t'F����B��IH��f�E*��P�[~�[����L���j1:7�s���J!cŎ�!xu�Tc�z� �i|q�\���x��H��R��{Z�=i��?����Dj���Y�k��'�a`ɷd���4�3��*���f%rζ����D|y\�����h�\��>?�U9���%��w��*b����"-DԢگ�˱������02QYD���q�*�ߥ,/a�oan�:[�4fx�w�A�L�~��=:��(��'�x��Km�w$����
����}�a�����?A`���5�p���̬�A]y��M��,_��?Q�o|�\
�&9�]�v��'}��r�h�l^�Sx���M���w	>�/ĝ�~�/�.�>�#3��3׷^�T3GK�\DI�1,��3���L����LWy����������:�F�ڙ�׫e���⓱p3�֙�h0o�J���u{��u�?��ӧ����põ3"��P�"�I��9V�����X�"7�!��e�1�Č`��=�(޺�[%�e�j�.��������@��"O҅�pjL623��nëuRVT(�ao25�'�ϫͿ�	�E����\�ʍ\!B��������Dd��MF�SX��lt���4��� �X�"��k������`��>�Y�×�7�u�6��l�d�ʆ0:!��5�%�o�af��5�KH"	t]�P��J�7b�C��t������?W����Ubal�{])���N�;�����Q�nw�	�K�Gz���t��JG%C�>�a�$b�Ƨ+�]0�K״���a�)}O
�U\�}�?�B�v1�Qא�g}~�����N��eڝ��=~�й���dn�E{|ϔ�A#���<��(!Hrc_�Y�E�q�e�Kk%=,S�tQK �r���g�i���%���}*��讝L���T��&T(%����E�0AZZ�ȸ��#�=@�R�%ߒj<փ0���k�����^��T�ֶ\|����DmH[�Ho�\�`$�AkB���X�	���Il�j�ɰ�E�����.�)�m�Ei�,R�Wˑ����<I	{\���� 8�=��9~U6�;E�g���m�cK�% %��RDӎ�?���A[]!N����'��x�����|p���)g��B-dT�R�_�������ٜwQ����X҄��Nl�C�:_�M�@e/�<����é��*�_�ag/kF�Ø(�R`�����<c|�4��P�coljܼ�	x�/f��#��뼳7����0�|�˗9i�5N0\c�����E]���N ��J���@|m���+��
5�6���a��*���M�_ʌf�s�<�Cy�yVڏ �Wq��^=t�V���S���GP8��?���ܨ�IZ���дE1\;�2��?��8`��&���	o.u�kYw��ٸt��/8r�2����;�ѐ�^����� A��5�(��pcK��Xz�m�2���#�@�u"ݳ�p��v���9���K����e](/��Μ�J�(�C���ob��U���ɤw�>f8^�¼��_v%��{\H�����t�q��UU���*vUf������G���.=����6����C�B��l�ψ����ܸ ^U�Z_4��^o�U�*�I���u���<Q]3:Х:���`u���y+�䠵�dجN�Ӄ`k��n����NU5�6OgUU(E�h1�����is�~�2b3:�m�����P�Ŕ#�k*G0��y{�]p�RӾ�kp�d��t줸��|���D�6tsQ�z�@44��l��5��c[�nE�i�#CC�&C��TJ>i�@ݾkmY������Z���l�6��!#&�4�r�k;Bk8�S��r)g���M�c!�~��:&�/�����:�l�g��E�Vf�!q���DU�+�ak�E� c�(��� ��7v�_��ʽ)�����V�v�_�[��K��.�!�y��t|�������ɐ1{��ljk�5�]��R�Ʋ�6���`�B|�"��M`���#������?�BLք�c�B�
EhLLL$�]+�)&�fj.�UÀ��	iWl�Uf:?3���������G�6�oz�ξ��̋l�Uװ�j?=.���K-ut�r�,�<<Z�d]j�4�oi�W�_�gY�种-����#"R	�8b:_���.`�,��I���:U�$Vbf�0����sD���z"��Q�ݖ?GF"o�=�c��zX�)?z#��3H]lT��^#P(� ��D�AҞ�9��̄"�	����N�� �q�>a���-���zڄj���P�ӕ%VsV_�F/ut��[��\{�.`�fq���3��!�2]���á����n'�~��'@��A�p5Sʼ�p s��.��Ffa��'E��>Kz��o�p6���[�&��9��Q�!�~hq�䬚�n�$�Du����u�j���sO��b[�>꧒uͽO�H6� ��@߹g��γ��޹���|/I;J���xb�J�Wʄ$ّD���Ӳ���@��"��6����$����jZ�)��Z~���KWI��_m�o�P2�-ɜLl�����Ư��l�g5�+H�	��ф�c����}�o��~�۶�{x�5?�0
�/9#��ѹa�95���Ĭ�$\���`$�h�M����B�_�4�ض�L���-�;��_�|j��ÿ6|ξ=-�!�5*j0y<���mN�dkk�/��<��Ff����8ǋ��EE�P�
�sY��nmpP?���&�~x���d��$��{���P�
2�'@��@H8-.��Ǔ�IF�f��/���2[+5���13X5�{�W��d�����U����С1�ݤ���w8��(*���HkyKJ��]g=f&�1��<���# �ƅ���H� �\���ݯ�[�"�7��&�B��h�_,U�,>Υ���+	ݔ(>ߩ��˚�ϳ�PÎ_���������l��ۄ������X�Z�f�����$�@S��Ed��k{�rT�"��h���������~�U���Ч��W~�#Z��������G�L�y�Wz%
�a7�y��4Rr�kVQ���5�C� �R�����*8~hʬ�K��aX�0�@�$[�����^�Zf�d�!���<1�]����ak6��Af�4��;��i݆���AH������m�/�Q�&��ǵ�-#EM�
����1�$��\���Qu���{��]�&�FR�����̈�����'�c��c�����*2���'��+���N_K�U�V �wM3��?��sI��S�ڽt�6�"�j��u��]IO�+V�Z˸�]W@�s僓����ƍ�����톕���0��| o\�r�c�Bheߩ��G&8����l���p����l'?�����D��P�ݼ�����}����b��-D���]O�&PF���x9׎��h,Z�',�'��a'��R�h���t�ꡋO�Q�ʨ���(�t���s�����1���3��%�#U�d�ʦ�,٬��S��+���Ӿ��"���hv����'~�]��3]����u6qɈnnP�����^���I
*5'�Ϙx
RF.2�� {�䔱;L�x\�R�F��,�5�5+��EC�)�� @�)-��ߜ� I�iMñ�V^��C��#���[2�̐��)���~�k|����I�rD�W�i��k0�јc�B�����UzC����x{�����#������y_*'�+�d,��VHD�䒸3�ɲ�9ǐ�T{��G��G�t��	yU=��&r��$�⁷�X6���Q	��&c��\G��Kk�V΄���vU�`��'H��(;�Z�|���ve[֍�R&�E6R_t��r㵨�I(��� ��W�����>�C�5���!��7ݽ	�����7؊ulЇEK�����IQ����n�:�A����P� �g�����U[���U:�y��A���]����I	��}��mC%�N�y�l��-�T�kOh����e/�g��g�0%����g6����w:굉\c�H��~M�"./2���?a�qZq���r<W�v� ����&~�~ٹ���)l�R��Ũ��r1*1e�+�x�\�y��z�xZZ�nwr��֞�O�gK�;t�f�W��-09���y���o�2��A�5�f�F�(z�c��Go<��AV�2�}�.031�<0��ux�z Bg�{O�b�q��_%k�s������k�FO�����{ ����4������C7�8\�M�\8�y��[ſ��^sMc\7��a;�b�`�{?����!���yj��295b�(.ߕ�ے+3���i����hiÜ��
,����6��g�B�^g�N?C�9�K���fͰK}T�q mZ�q'�2�΢�[��%�۠2R��|��G�q�Zk����)١���˔�Xb���QYS���.Z?��C�pu�*���|����Qif'ۧa'�����!"�6��tq��y-���m�p�NloNO2ś|��Գ0@�I���y�	�\n���dg[�� =�������E�����VU��AN'�1�!�Q1nZ{��f��kGF�z�����z�K�;����V���G��h9�����:��$�ۨ��|;r�L��n��N��;��Pܖ/�-��u_��b��E~��,7�$��mSm[UEx-��r�\$nk�zC�ig	�������ʮ��!I._��i�sc}X�\D��9�h�s�	����Y���D��g<���6�����>n�w�!�0�/��C��6��`��*����iE��7pa�������z�z��R��?��QlT]�#���ؼE%�C�LH1p- @�w���}.mEc[+��&6A�H�Ϧ�d��*�0(���r���y�V�e`�B2I:+�m</���|�<��Q�'AS҇�����ZӆX�6��t�d�14EY7���[W �el	�/�k�����3��^Z3���*a}�9�����vnX�sF���n���4���ke��ȸ�{z��Ò��/��2u�u����e��Yl�|X������`/��)'N��,��
��*J����@���X��j�a���$C(@��S&rw
=d&��׆5i�@�ݛr���9p}��k�˕D���´x
�/3 �|��?qZ�"%<��P�C����- ��;�ֲZ�^	M���Z\�s���+�����l�7R�7�o��L�����V5�w1��Nw��`ʱ���xDȯ�KhQ>�c�9N'�9h�Z��I}��+鈩��-����|��0=&]��ש����B[[t�Q�[ɦp�8���o��d8���Yp�"�/ͼ���6w���Rέ;��Qp��?�$,8�_���cM��Ce7,Q�w'A��[��8���%2�1"f�g�ׁA�DH�����W۸1������+���,@|r�	���é;�fQ�<��E#�b.8d�Jb���?mw�7�3�iJ�U�ű�ڵ�hzgG�<���q���ۮ�ǧ��煹\�U*0�<�퐍Y�V|�;o����MSЀ �ƬK7�������ud}�@���*^v@�l���.	�g����6+��	u�L�G%���އ�y�DϮ���L-;��wvֻ��E��Z"P����4o����낡?�STߘ2˩��N�x�OK �'*@����s��|�5���}ub��޼5V��A��^��������ٕ�A�Ea�z7v����l���$�3�,����+����[?=�X��}=�Il���x��	�=�@.�����+�,�lF�	���j��yR�DW�Qz=!D�,�QVׂ�)��ϔqf��4��k�}��D�f�\E�aw_P(�5��O���5�ɱm��9��E'?ɬ�1�M���,�?U�����k@����k޹�[���O���{��~G�ˮ?�?����2���٘eLd�L���m��hwݨ+��MIǼ�*���U��x��?YI��3=��s��d3�dƾ�$?ʳ���	���G)+�=yT��b�rfMt�>D
Y��Y���dֳ�+"#h�n	�"B�}m+�/{����n#.�(Q�kx[���2� �Z��D�J��^���1��p�E���<0Ս߯,s s�7<$�!*��C�h�7	�mg�`�s���6Ƣ���\�^��%�*�v���$϶Y/��v��U$��l�1�LE[[�t����}�]�°�ѡ��p�����z|�G�����D��;շ��ǔɂ>���8�����3��l@$I\�|���-�*8���z!B}r%���hR��'v���2?�w�N�B�`��M�@^x]���������Ъ�m;�`�Y�z4'MR�.�9m�-�cP�����N ��I���in�c(��{������u�� y�m�i�Q���q�;65?}JC�Ix}۟��l:ii�\�?iuK��S������y�]���b����KR��	�<����u�!����;"��l���&8�&��s���߲�a��$WE.��q�e���+�>�>���m��!K���yJ�_(m�?�殒<µ�E��ߩe�>��{�K�80@e���u�|!�U\�>砟f��2+܀O���T^��1q�Zy������?MK1A2�2RTŪ��5Ƅ�����z�-��n�t~��Wcn��i���q���7��B*��z�`k[u��Z�l���1�я�NN��5������mT%�ų�uئ�%�P��CB�ZVC�d��H��f? '(^�|��?�53��6lC|��[�m�'�q����ݥk�vz%�6]��S�"��%7ۀ�]�D�fX���g)�_�N"�	���j�:�{|�4b�}b��g�M=d=a��Jn^��\���
ӧl�ךc�3��R�A%���ಭ�2�ř�X���a�f/5IuG��Eț�=qWKBW�������1�E����g}+�飐������/�0I�S��+�M���$�>�;��)B���ў �6Z���N莮*i�V��w�p�7Y��#�c�B��{q5r�d�v:�!֊ֳZ'{)�o�m�'�S�wh��,��������^���������[Fw��F��>����`߬O��ѾR��6�E6���t�7}�e=֟;��̛����� ��Kޝ +I�����3��g
H__�2��E��'?֩)�y�$ˬ�N�'͆6��y�?@TU���z�MV�������}<{�J���xё�L7���1)>���֓8���������gR2e�}�F\0���C�ۉ��ub_�b��3�ꫩ�PzQ��M�h����تX�K���l���~��/�jh��d�b���A�M��Ċ���<t���*.���O�ur2�p�[���=�Zu����_���i]y �G�GmLv^[���Ҡ���u�_��]y�K���ʤ�fˇ�Fap7������h�`���Jq�f�O\o�I���8z�\dU�hs  �#IkD���O"���m��M����^�	3Y�s����,���<4H�J좧@5f/�������L3}g��)�!ؔ����yP�J�u|�}��q��&f��ZG6vΣ��EHֻͨ�v=Sr@�'�uȉh'�]���6�i
�K�33
U����̳,�+��(���v��ԫES���ӱp;S؃TV!��5<���m2��\�T<ev�Xl��{V��Xs�I�z/V�-�'~����`�xF���1\��-�M��A2e�͓�z�Uט�j� �J��r쑵�����}�\����+�!�p��!K��G��j�t�J^�DM�{��f`���%I�6�?\�Q{�C�I(CA�-����n��ݞﴴQ��Kc�W)������$��+��&��d��2�M���s�H�>9�\W��F.�eM�y��5�&C<X�⽶FqY�y�+(�[��/l���Xh� f*i����K���֨�����g0����-�H��d�I#�m76�X1�~*򜁽=����>��I���q�w�:/mh��82F���l�%=��v��Qȵ��jی�F�挹Y�y8q%MLB�k�X��RX-|������e��4�HE~�`8y��_�C5��T@��\�s�]zׂ��_��}�$�Ev[���5����c�>�/�Ưڗ�{��V��`J�@>g�������.���T��v�X�M*���=�<��
��,��l:4�Q%oEd��ig�X��P�-�[3�zQV�]��^�Gѱ`?�>������}݃�1F�u��!+�s��S��1׿�<p����]��k2�Ev;��qs�]S�:X��㺯0[�7�¨g����Ķ	`@*0ڨh{q�k>A�+Zpn��ύ�Z��o���_�<�7"��7��!3��iB0�b��:����������L�x����O=܌��M[I�d	�G�`j�ǃ Ǘ#;S�,���m�D���o��ZS\�j-��
!�5p�[5.��<��'���}����<��w�:����� �8��9�.�[��ǻ���3AzoY��.�~{bk2"���m���!5Y\2�d+�K[�^���A��y� &,�f������?��b���E�=(P<M��FvPr�z9ӻ��I��t�>o�j=A{6��eJ�V��a}G�|Q�T�ܺu��;��|�Z�}��X����a��G��/�ME�tj�W��Å��HcP����v�ȥ\&7#@2���+-e��xm�D�'+������˚k���G����Mt������{�<�W �� z���]6�����q�Q֊��fQ�v3��������:����ĩ�B�M�h�@f�}�Rƨ���6���]秧"�q�zvȮ#��v��҅��S���2u�����ۆ�9Rd}Y|���'�����f�ua���V��@��x�j��|��]Gc̎W򥐢���;`*Q��h��x=ȅ�Q�d�C�C�h�W�׸lB�'�c�v#�/�e,�����&�!�d���w �ǭ.X���lT��8"��$��i����/����`��⧵��5	�ѽ�8�Cؠ,�0I���luek������;.�$.����Md���I��Q*�c�.$-]�	�=O�o�-�K�>������O%_ZM cc�塮²+�G�(�NGpT��d(s�6��ۨd4f�M�W�%\�OX'�j��^Q�1q!I@��Z(��DD����;$��[�S���.�ƙ���L�	��lg�2�D�S��M���͗F��Sئ����B2�1jz�"#�].�b��]���k��1i-�!�ˋ)�8�|���Y�Z!Oѿ����F��q��F����V��7�<w{y�<�eE��c�K�NZ����9�.̨a���
���)��)ٸþ_�F�07�989af�2��"����.��w�n��a�י�h�`��� 
Jw}d'a��;�����_�-�ϲUWu�����8�E ^�E�HA�����|�{�^~hA����&�?������9�C+ab\l~ڱ���'��n]7h+v�l�V%�5�WbO�檔x�#�8�ځXS��Ey^2�9��) ��.]��( �|<�o��_���h��9�����d�7jA_aFe�P�N��E,�H<b
 顶�:%���a?������\Ѓ�Q5�#�ow�=qW���5��I���`c���[�`�-�[���ܪg1�ۆ�jDb�P��cW�Fa&��J�:�t,9c��^�I�Խ����/�4M�؏��C�3%���P���%����sAD�s��ң�|�c����N����F+��!ƴ^��M�&�ϒS{����6F�s�ک,�<3�b�s�T5@*���m�J��_�p�w���#��v������� ��v,�Ȧ� ➩�N�sKKK<���Qc���V;��E J67R��Ւ�w�'��'�8Q'�k	��Ł�A�د���+��o���\�0N(�āvw�R��joK%{E����`>I��B��?���ĉ4s���V]��6=,ܼ�5-,:�.�덺êY�"38P���ę�i�g�>l���d~�A�F	�*�_�՚GJOk�Y�p!?V�������v�<�@g\8��X��u�#�LK	\�U�n^TQG�����M��XN�m܇�����7#s�w��1=��\HL��q���/z56�� �}+1�����ͨ�k��EK�Z�U�ks��7��D�vk�~v����tcI�]΋�ę�����z��5�u�2��1ȔO4�����Q���tQ���:ڃ��P���]��i��B���gyO��xx�-���Ӟݑܶ��/��y)f/���M�o�
 _��}u�E:8ZCzf�2��[��U�-5�|ZW1�x���x���L�%��:�T��M��8O�ͬQN|�R
y<�b'9l�%|nV�8����ꈌt������j�	Ŏ>n��%��
�וG���Vv�5"�㫄BݔUv��I�e8��c�g�4q}�����ݭ�p��� �l�Qm���X�w�u�_ɬ |p��D���
*��yAt�p�)Ȗ򽍖E�P����
�m���4D����D���0 |�^v��ōq�����YTP�0O��f�е���8�H3|L��M;���0���̉и�Ö��8ω1���{�ݰv36W�W�3�70��lM�1��	����9�r�l0i���_�������tGv�����5��|��K|�xK���j��i�_�of�9���W���|����W,�T�ot$�`E�%J�eTR$�j	v�C^sd��"ˣ�4]��t�Q/~y�4���d6��u�����
%O�\xPF'Z����Vh��f�ź0���#a,�!k%�����	��"I�E>�e6n�!��e[f�l�P�BQۗ�mr�0�����.���D����P��1��6���ӥ�>4�s�����c�7���p\fEޚ#]CU��|R�eU���P8Nf��3S�!��</�H��i�@ę�L�*µ2���0j=Jsm��e��}�d�:!�����XI0{�4{�G��� ���h�א��Wˣ�E�ބ�53���/��n	�}Ԧ���z��2�#~��5�_��_4/��L�TߤB�̿�o)���U1A�5�5���J��*���te'���$��v�%O�k��`���q�[��O�7Bs,���Q��9����R��c`"���Q��0�����Z�s�%|�G���ɽ�ŝ��x)Wt�L�n���g@���ʕ.����aHC�2#un}z_E���9��������m�y)M;]?~Eݮ�UȞ'��g�E���isQ���`к���Ź�Ҝ ��=6�<�@|�����D����S�u�=��7x����S451U�7<֐_"�g�o�θ0{i���wr�	��?�{��`��5����4�I<��uU����)��;�c����KMh�m�څ��O��~X����t�X���r���f�=�v��걜�
]�A}�:�g��	�,�l{k�m�	�;u�Ӕ��&l�B�*]��9��Fr��O?���@Ȑ��'�vsH���b����͏�<I�[t�'��$��?�/,&��|��L��-@*��<`^�J/7M�lj����׌��F��1��3�
F<}��E�i�Km2����!����/�'Ve�}g�*)��N�p`M�P�Nw*v�9��rߐ>�J�^�+�e��D�dnػf|�ѿuuR�����N��P��hj�a;�&�Da0��	� ���!�߈}J m=j9�*���� pH ��0 ��$��4&ЫM�s��j�ɩ%�J�<�h��yv{T���

9`%q�X�8�׏�z+�d������T9�g������Q�!ȥ|����� ����b�c'���@�����4�"��O3��c�}���V�c�솪��ݵ&k���t���ʕײ�6
`�Y��G=�D��r����\%b1Q2e�S~�t0�?%9�������1��set=� (~��_�֯��������U�����mB[���\�em3G��g����kD�*�7�ض���WHܼ����mt�JA7.|�lg?�:b|��.pi����ޘ:��Dt��L���YHA���j���S���:�K+18�Z)��Ƹ�G�	��<n��0 ��GX6���]��j�I��h:�N������i-�;n�b����[Zo50�.��i�Z��d޸YJQ{0?��@J��眳��oX���Gb�̻+�i=2c�<�bl	~�nZ>˜���/呓kN����!�����%�dM�U�-;oꟾL䝈j�kXhz�)�h��	�K-)���B�^k܎���ڕ=���1C)��1;%����j��1mc�����7ۉR焌�a!���V}��N�����ԣ9[x��&&���g�7[{D�O��9S�A�/�NS���5'��n����߃�s,�m|��K-��y�׾ѵ?T�j���;ZL�ĳ�Zw�DO��o�g'|����(��:I�d�F,F�M 03�d�ը�Q�:(
���Z�ܶ���]З�=�r#6�_8���O�7#7I>�����{��Bg�:��*ڥ��3~��q���-�4<ɦgj��BF0/���DD܌�>D,&|�M��dܭd�kϚ�9r^�S�b��Md{�;r2�q�~b0"���L��ż��#�|��$?�*�]�}���5�A/1���A`��-ֵ9�ic�����~^/��� ��lߣ��~-���b�4�x���ߴѦԊ>%�����>yyl|5�ڿ��〦d�/��9��ol�������!���h��������z";��%ɋ��	��h�и�ɶ�@d`�f�H:�ʎ杛�/z�匵Ps���E �5�>˾��qd���'X*�&l�P���gA�uP�j%�}��i�cVm� +����Y2���W9�f��)&�5$w߷�ƓF�MR� �>�E�"�_7fÇN�Z�ᨓ��!�9�J���Í�]6������>>�_Tm3n�\�KE��%�u+�C�A�kF�t5ab1w��#�z�Z���-璇o̺d��E�<,�ު��>YӾy���#�փF���+
N���e���{6�[��ǖ���A3OOʋL��`9VB��a��	4��L���ȚY������j��]Vr�sXm�<X&�+�Da�Ku[�ȏQ�r��!��8p.�x�V�|x�k�;"���PM�xn8�g���5G,����P�'��ҧ��_����'c�PF�)/dHaBi.W�%�H�������}&3�.:�*#��"�7�#���du�;^��p��J��6�ب!~1�1�	:�A4����+⳼�U��Bu����w Ǽaf����[��M�Da�߭zS�FP'2�3=�����fk(��&��>��8�g"�3e�c�D8rh��@�u��o��^�H����'�}������ߨ%�&��#dl�nz�p��(�c)Ȓ�OH?C�?�}�cv���*�}��J�:�4�o6�
p��0���6��j�3=�I:Q"�d"�;9�	[��&5c�h×I��d�������_�)D1��tn����p����#6ב��#6J�.Ef{Д�W'�Թ㾐x�αt�Y��?�X�S4]w�C�dcyS�Ƨ,\녍����R߽�`�rX;�.����Tǡ�(-�јH0�lBsp�3E�H��l-5Ń������ŷ��;�P�k�0�Zb��oYxlc=�ސ����@u^�ކ	���Nm�ír:rM�W�i��mb*͆���$��8CTVP^6M��DD�q-%��ᇸ�%{�|0�
��JzΗ�*S�C��6�������o[8���D��v�U���+�~�s���D���˞��Pz��Nj��D�#��D���Fm�K�KR �eҾ������8D��:/#�� LǤ�)���1��Ѹ��K�|^CaUnF�<�k�i(#�9��fY�5������UZu l��܀�_1@v^j�y!%}Id�r��jo���*�Ӏ��/�X5Dsu�O|A$C'e�m'�����KLL?䞾�$�Z�v-֪����M��c{��U�w��x�������E����8֦3R乬���H�>�b-�vq��{��𰤵�Ұ�d� �� �^�6u�۷�b�i�j!�po�i��J�)�?���b�j�Kڸɏ��q�#�*�X��t,#�|SD�_o��RA�7{?��Y�q� N
s�������Y����|��a��rV�(#��%W��۱iJT�u@Ԅ1��!ÖY.��/�:X��1����(>����6�C��@��+d��Z�{G̞��)�l&����y{��n�֫k��46�f���y}�.�.�㔻���.�*����FE!��5uz;���j������O�����������}n,:'��$���T�'������/������@���5&฀�Y_H��h�	���yG[����^�������챪.�:�� ¦���`���9�ܴ���j���L�H�O��?� �d���3P]ґ��(�@X��DW$J��
Р�9O}N�C��\F��s1�ka�S����	����Z����t��
;�i]�W���E��H$��XP5�"�.��쿀����SA�m���rƚ־p��u�(}�٣�ʨ���@��I�:lL��.��d2F9`(q�y|��I��6S�5S��pU�y��8႒VR,�A�O:V�BЁ��36p�Q(��h<���|e�͒?�3x� ��D�]����
�f�񾿯��Hj���X�v��@��!�]^�ՓѱaI@�űvC���}��7���7�:=u�Y�r���R���ڈU,5d���wc��V4��R���x���/���%Fg�p&�iE�������FŦ�0���<D�\{j��y+�`�8�}d#�R`�ѭƉt��ou�0�7���n���XFbդυ�ιD6�Av�L+�:0lj���1k���s����������� m������w����m��/�Zw�ꠧ9+΅LGqu��JF6�x�u��b��cGB���:��eM�Q�7�+Ղ��8��ꟃ�'���[�>v�V�;�{�}�q��r�%jω��zo���@��j�ypy��O[x�u��3B��,��	���$"O�).}�5��?J��9I�f[r���q�vG1#�U�l��EZ?���F~�6�t�myT	ߣ�i�d�6b[#�vj�rq�u��D�:�.�&�~�\��X��*�v�z�Z۷�w�>����$T"x�*��e��

5���ꭳZ;�}�>� s\�v�4�C�s
����I�'��$�{���6��N���K�ξS�@/쁿kHׅ�
�Tnic�Ⱦۋ��ja��x��k�'��W\L��nt��Y�0�N�Э���'J�[�x5�0��N㯉ϱ��U�	����$8Sd�v�&g�t\ݙ��5���!�o58"5c���8��p��;,�-`�f3���t�Q���'J�ӱ?�P�]Н9x4���Y�0��!����m��˗�G`�~_{{;Sw���_�m[a�g�?n5���pt���N6*���8���Q��s!�"ڸ���sv����߽޽5E��?��1A��RB�~� ��?\�<m���k����1PH��u�a�׊���I|�zt�sE�$$�Ԝ�m�=�⯗�ɓvl}��"�;C�燇^��X��#Og2?	�9�b]l_mm��/d���	�`��������`pg1�ia�j��ݒ��Rk�g�[��#��߂�zF!��|�?�XO�¥�Q�;~�:��cg�t�^W�/SD���a�OJ���Hî��0��K�k+����CK��!��L���)��-�D����3y��B���Bo [���3��3�s�E QS����
�+��^�8����}�8�D:io��DPWk��ˆ�M�����N���5� �fe��k�i�Zu{i�T�F�i	�p~�-H��֍�n�d|)|�++M���8к�uj_Z�蜐�ؾ�<^h�07WK��-�{$H=�9 �S����Gf�,/���/��/�*�4Y{��o$�%7���:v��.9�9|t��,�2=��	!}�ϗ5�W$p��T-Io��s�' �����H'������Vz��:��]�YB�RLPs��{Y��Z�K�l�xѓ6�b E�U���´r�nv�B�M�������� �4�}3���Q���-��*pK�j��X����h� ��CE�!���v���쥓p�|9����c�7���]����|9__ш���Z�ɼ(��B71��)Kd"� �<>�i4�Ńx�4��+_��yeuӱP�����-N��,,���y@�B5��I^��뼼D��W� �V8�ZV�Y?W��	H=�'9c�,�8��}S��;J�=_$zsEU��M��)�"1�B��|�B7�Г�6���cF���,�/�����n1�N'��r����#|�sCc㍪j��?����z�p�($��'��e��'���bMB�����yS]�|׶Lt
�)��4�o�)@�ϨΌ�`:���	�>�bNN[$�i�;����2܁v�0�t��6YW��v�xwe����R(��6H�X�(@|s�T$[9a���D�X��DW�����;+
>������|�5�N��K��D��N��f�V������-sB�K��U�'�!=�!<H�hp|J��i�@���g��1��6V]�W|J(�k�x�o��5AR��'+Vǅ���O2���̦�ǂz�9�sn<4�` nK�q����J\��g�o����'(�(:`������A�et��x�Q��AX���g���J.>�ܝ�c�#I�Lt���oQ�~���2���/0�E!*{��9�Jٹ�}w��|�4fF<j�чsMȲ��%k�8tv��"����<$J��
j����ڨB8OR��W.�$��=(^���������?h�y���
MZ{�q5X�g[-�Z;S:�b�TƷ�h�͆��vy���p��"��>裿嘕�>=N�	s �8ʴ�� zI�b�7X�֔��mU5!���X�8}C5����P�p�8h������s�ryh��z����Eu�ض�tun�y8����~Lu��)aD�R��%��ߝ^����IlQఽ�^�
x%wgZ�2��TV��򮧩Zw������eD�c��tŢ�ۉz)���|��O�ډX����g�n��!od3Ȏ8}F����������Z�28	U�:�'~�[��$�@a���<� ��[�v��L�ErI/�OY�,�\�3�C�$���RW��Yx�AN4(V+/tm���r!��|S��G��(�J6V�1K<W�Nrk��s���ˇ*�x)	tT�Nf�h�h��/�=�5��,�j�u���"ݓ}��Iyv��mVt4vМ��;=�}yL�=�4�N���
��hK�:�O���w[�g���Z<�W��hş'�z�<vR'����[��f �D���c��y�нa2Y��y�����.t�!a�.a]���Hz�΢C�����#hh�W�yoK&�����������&�=�JSC���O���=�ޯ��8[�1��0�g ��KE�,ɒb}C�kY���`��󉐆8�-��r��>�F"�=��9�5�,u'�hV����r�1�Ց�f����D�݇s��KVH��l��~����2Y�E�.e��[�n��Z-���ȡ��Ķ~����Ùq (�F�K���g�-+sR� n#�Һ#��[-~��Vi�_q'�U���8�|���� ?b�;V"$Ɛ�v��_��E��)EETg䤿њ�1�H���@� ����K7vPCzml�h6���4[q!|��r�x�K����[��U��EuY��d��~k��+�Li�:������½��:��ݷ��S��4p(�j��ͮ�ˉ�q���&��f�|�<��?�m����[���*b��c���}�qDȘ��'�؈h��h�Ϯ�{��>)o��L��s�����W�+f�ur��CĚ�[:z?F"֥<���Lla����纥������^�[���tr]u~Wvh����E� �����8_���nn6rv������i�|%���יM��Gx�m�?9�N��qW�_� �Lwa����	D'����n�&�{�/�C���7��"���Z}������JU{�S>Y�A��J�\V�E�o����Z�����~�K�Y&����B�H4peB4[�f���zZ���aX����滦Z���e���g�,��c���J�gZZ6�ZǤ��'T���/	�
��V,�QdQa&��zݙ�ӌ`�����k�R�W1n N:!Yt� E����y:�'ldp�Pe>���;�~�j
+�En���������Յˮ6�M�<�bN͕:����i��F+b��6��]���&���qK���Z���f��f �;�����=�ԙW�A��j�tne)��o��!x멉�ND�륦[�4Z�LF�~Y�Z���
�(�\�2��������W�.����{��?%	�ql�l�LϬC"3Wo�n�XĜ�b27�i�ˈ5^@k���`����E/�վ�҆�`ݠ��y�#�.؄B���z��;�ѿ�q �4�Ɣ:�m�~n`R!d�g	g�\L6�9(�T�pKgz>�"���f��u�D����WnSG�o>�&��}��$)�>T&�H�������sQd�# \��x���\���%DK�$J�~8S��-|���j���0ۜ�zqC�ko�⏬c80}��A1��dO�n�X/`N�<�@_]�y5pX�鯗zU���/7�4@8뫂Y�2p�jJ1�5Rb��#��_���`O��>�c��@��� ���'!8~�{u�c�����@��!�����,����]K���u��_����}D�N��:�:MQ1v	���ꥺi��w�t��S�3�G�͉`�>wA�o\��7���/V}1���>�#�&�Zbh{�يk�dS�Q4]�i���J5Bqc�������[E�J���(x}����r,N�����l#�����V�с.�4��0��aS�G:4!�yjd�y��c PD�m�����UURu�i�=���>V�9r�Up�QT��&l�ّ2_�֍�%�������DV�����/����=����ȴʶ��k�mU"-\�<��r5�)s$9�İ`�`��$�R�Dӆ�,��G�M���Kf`Y�y�b\��v�6�5��>M�R1������k6⨝��-�,h(��@��\DW\-�[#>��ƥ�Ӊ�� n[�?�6��#B3��w��9�hK_֫p8U�z�jeA��F���l�(����ﶾ�">�+�;�j�4[÷L�u��V�Yfq�9�os���J9\��b�F�4v��cw$+B͑���s&4���	T���&��9D��i�Ə
���Q��"zD��u�S��5�4e���h��-�Ԫ���L�(�d�6@��Qt��nk��LI�2�Oq�v�is�pR�c��)������̗F.�`�n/ �$Ͽ��6jI#首�%�(�����s�*x�g+�KJ؜��"<n��Vڲ	_Sǉ��	��Z�xOd���Z&˳������˛����_��7��v�����ʸq�CN��Ӌn�ҕ"__�O�D7�UA��D�m��z	�&:�lw6�"�X��J
�֞�u��m��o��#�=�wgm�$�e�ν��X�0u�����{�?���'e�)TOԸ8]�h�7�����i�=_�~Ik���i�A�;��.WGޠ�������@��ם'J��:D��TΠut�)�?���G�~Ԛ��'��?E��O0	0�� +��l��$S���i/��fݹ�%>c3�W�eg5�� Ӎʄ?�`��r�$� ��~$��_n���U��M$�,��ĘW©Gs�\B�<����~�NBM;� i���D�{�_��|*�?�]9F��{>�JY���(�j�9Z@��Y��Ӵ~j�3���7{C]�Wp8��n��c=ӐA3���!<����#X��	ҥEF=�	(<�M	�2mYu�v��G� ����qq"VP��)�y4]���e��Hܝ��F^��Y�Ls����7��H�Pz��d�!��6�8��9���	�D)�պ��DhY>g	�����5���<_�[�Z�ۺ��c����Ǚ-��I�@�*�,����tm�+R?�`�*��_�M��Μ_���z,����R�o���g�kNݜ�0L�"@����7���4��bp$�o��7ࡓ(���u	"t9c�.`�\��m��x}E��AV'�o��@ɖD��.rhw{_�>����:~[���ޭ��'�N���� fx���K��C�9S�t5�	�986����N��p{�k���>?[�����I�<��&[��@B��:Y]��m��3�Xm�aH����O��"�Mƙ�׷���o�XU�� �� .����!���ormgZ�˼ӆ�C�<�z�ς�[IR���ŮD9m�^� ���B�Qk�H�+"!�9I�v�ʆF&�34~r����>���"��qi�
Ur0������78��t�'ޛ�5�O������fJ�C�=f	O���y�;�mطVǭ-�.n�Y3EQ�J�����(�G�
EQ�Ĩ{�E��U3�Z"v*�B�뾟�=������<��u���\��s^W볃���?E�ڍ��ϰ-vt|n~64Ky1~����=���\��+���{<}���d��褝�m�.`�I�<??~�Iמ��g"��݆_����ܔ�OPW{�g�k��Hw��|�1����t�=�\�3O���|7?�~�b�#>������e11�����q���|{%�esv��'N&�~1Z����C����8���a��x��[h�� ��`�����y\�A �n{�@������y��pz����J��]wi�sqw���*�ֱ�]]~x�F���l��4ݭÑ��	��Jd��˯Q�M[cܿ�l�t��x��w���?�A�)ײBb?��N�����%3����������L-QtH�[57�Bou�e�ҮC#^�Pft�8�;Wu�̢�+����S�Li6JF���\�W�<#����ƍ�J������VA���¤I=p
q?�� XFu(D�ha&Y�Ύ���?���G^-x���]�s���+A������y� %jMo����l�Z۟J��mї�¿�zM�uW�-$,p�W�������uƄ42D�{lu-��^������� �a+�J�敷+�on^3P�N�F��P<�p��֭R�yY�(�ӵ�ކ� ��タw� )3�'^��dIV��K?��� �-ԄZ�&S����y�#�Ʋq��w��|�B�.Ww�,��E0ʲXq�K��Cr��p�m�V��l�#���J1X$��ߏ-	T��/�>deo��jEm~ݻs���CF綣�����S��bT�9%s��,���+�X������9�0��<����t.^�z^H��2�^G���>o]Cx=T)G���lδ� ��.�X��m���}�ЂKd����@�+Q$3(�a�h)�=:�k�돝�eΥ��GK����������~w�@v���4�bEL;�5�@�g��=�#�����6��s'_s���χDS�,'�Z�'��+'��Q��y�G�c�[b���M].�&ڲF��s�O���?D��j��{�{�_��r9�3�U]��X�m�'�aq2'rzzm�RG�����-	�3�%�Az|�=�B8K�KX�gaz�V�>�7 [hڕa��3���S-��C�J����ٮ���k{�h"?��w�mrQ���Al�f�f�j����Iw���_�U�-¹�
����'�0��\�N��"fh��!|��r��4����N����2vF�w���)�J)���Ign��F����i�oV4fǨU������qV��/  w7��|G��%b�}��LC�V�۟�,��M���}�M��k��v��v���	��gE
��-Z'Cx$9޺�n�&�=Gю���hD�j�m���:��v�fUĬ�	�ȇl�9����OOB������*}�ښk����=�vM88��O���Prε���FC��'�΢ƅ"+�0������+�3��-��╛�/�sߝ+C&�v�^��}���K��o֪yp��C<q?���H���O�{�|�1������rB栰����"y��4���2�@���e��g�����棊��*&5�����r�Α�%~An�}A�xć;��nLI{�  ��|X�(�V������e�y�&�l�����x�NWPǀ������/LP�{M+�S1r%�pM��L�Zk�����u�g3�r���h�wuu�r(�;���5�a@T]��5g������"���	��\��,}LC�����㉠�{�˞��.����r!��$���a���SN�?�������Tq�wb"��uTK�H|�uɌ��x��ZLY�8w��A�LҎ��5PȈ"ȖZ&H�Zz���l�1{��5*��ci�Ӈ��(����ǫ�(HN>,�!:��]~Z5�f	�c1����_/���n�2Ak��#�}����9ٴځ֣ *;'���A���+����:�@q�j�/�8xG۵l,�O� �+�2�����P7��%��t�"��v�5�o�&*�IR�g=�p)�� o­����44�:&����2��&;�<��������_�β+���L�P#6�Tʐ�sll�Ǵ�����"5�^o�5�vyʴx�9<)	=Ni﷠��l��ݹ"�m�=�RcH{�|O��E�ǲ���7�w�k�е՚;L��?��,�	���;��h��7����@����
��6����O��8�p�%��d�<7DP1�B��3�/�s?�����f�����z���V�~?�j�L �9�h�����4*�b�lD�D����+\�_���Q�؉���JJW�$�m�O}~��?j`��6�����0ϤK44B�������!��Q���.-|�u�M?��?W@ Y��]_��Ө�f�U2~lW��D�R���a�5A唶��e_raN����X�PM�@��J�:8���7j�o���?��F���S�}BfF)��^/�v�:�9f�ڬ��J��,_KGW��$3���p\�t�D�2[�j�؞c��ˊ��a��q��u�#7dd����X1�Κzf���E�;��ۯ�a�9�	x����44O"sܦ���&0|j�̶�0�6�2�t�j�V�'}"�����NȆ��i����)�u�<�GJ)�Vt7u4�݉�5��"��X��9��T�p�"���K��)"��2ORS;um����hj�XH&��H߱��D��F{�O�%|-��{�����?�\1Lo �FJ�d�iM� ��(9�j��IIzK��g2�Fe?��º���͐�2n�#��dtL
�z]	�o�/2���@;�#���y��d����ww���ޮ���Rv��_�_����,_���_�Jny�L)2э���b��}����drcs5d�KL`?!�g�������f_�cS�5ŎR�Gz�榆��;i`0]�����a�bYT)�*e���N0���" SH7i�<h��N]�@���y�C��WHЦL��)?` 󚵵�Ƙ��R��#x�z`����	�����{���z�%ПK�&ˑ!��9�������q�})j��и	(�S=\��O�o�#]�@��*RԆ{���6��n�2Sm�#��w�9g��
E�}y�{��ـ�����-��6�z����ډ�nӐ��G"���[��1��N��b9��`� �h���jߠp?.�j`Ѿ���8�e�/ ���c..5)"�`٪;�
����;ܬ��̴܋O:(\�v�R�qه��Y�l��;>��s�IĵkBLn�a2��B�]�a��
Eğ�dZ�5i��.l��.Ɇ�w�N}�����qi�q����� �i3D�w2�j7�izS�s�����'���F�J�E�M*%�$�$�S��ٴ7�^�k��W���rZ���Rw{��V���?�iv4"& �E�b�Uo��w��4T"��g8� c]�>�z­;2��δ�L�&4�H�����ov6	x,��񭪸&��Ȯ���Jn���Ɨhk#�N2������&��[	V��r��Et����I���ؕT������k);�P���;ɼ,�!3��\�4Ř�~ߺ�+w������S�~̚AY��kۿ�u�(�c'��?I�_K�W|+�m�ʴuu6�#�!4{{}��wF)n�i@�0��Yt�ϊ\�L�P�ug��K4����uY3g��6^�#�0e���鴊��_�U��0C|��"�KA�=*�;C�_b�=��v�l��D�t�#��^q��p`�ݠ��Z�+.Z��#���)�dOKr[�[GP+�a�E��7�z��
�I�����H��GYX����k��v�W���k��� lf�rR������))K��xr�d���6W�j�-_S2�7*�z������뭞
���[q,H������h_dI�j��HL�<n����^��]~V00��I32@Z�M�m��0�E=yd�W7��R@hl�/�1i�TN/�$l���!�w>���#�G�x5%U���J���� ���w�������%��Y ���H��#���%^x��ʩ��s+?����~.�%O�a&!'`Gy>YZ�e�3�?)���O�z� �9���"��Z�D��3���xJ��N[��D�n�[�f&9�WҦp����������jΔ52���q��𚞪�;��/ɌN )�s��l�/fZ�B�� �:����1j�>���&��~φ�S�V�kC��2��W�taQ�n��Hy1!���p�����E ?_	�H����q<nE�.[����K*�e?C0������e���o��u��ÿ<NG_gh@}��
>�1{��SB�����*�����F�V�+��<��t~?��lT���l�����-��(�$Y+�\��ۤ�xG����ec�B)er���1��C�V>�N��VW�zO������5�\��ʉ4�*y�:k�'�+1Cǚ6��Y�b�I\�{'����@D����s)F�	ozx��7���ߛw�=F�5\���|���+m�Li:2`Sk�n�sj@��S�p�#�d�u�#�b�(l�>��<�s2P��4$(��nUt�z��xо^��D�����j��9*>H2�l��zakק1�9,lV����&�d| 9��"��3����H�~4g����	B��ٯ6�F�1�[���p���T4�����+{i�֯�7�߲��pg|���ڼ��_F1�B���u�&� ��T��0���~�V����7G�.)���I�L����z��fN�F�C�թ?G��� .-�ͼ��>q	$���l�I�G������ブ�����ѿ:9�k8+V��^�)Cm�];�Yҡ���/Tu�����i�N>i{H���i�]���X	x�`�n�h.�6CnP.�GO`IY�� ��et7T��$jt�Hו�/��7�1�ne�[�-�8�+�z���t�_���̩�T�}�nR��,��\M��1��(;�ĵ�=z�-�1�f9�دGH�HJ9�3�Ӊ�28��.�C����"e��vnss�|�;����̓?�x�,��uо6��`�x{][әK�}������6�P6�o�ڲ���B9i0[]�35N+H�/����jYZN�ϥ,�O6O;��y˫���ad<*W�B!5�_|�n׃�����������=�gD]Ŀ�����6�9Mn�ri���@؆gJHڄ���A-�~�=�ZZ�U3�!p+��HΧ�q����[n�[��ʔiB�F�������80�J��6`7d=�Dg8����,T"M�����Yqk���ͩHj��qVخ0��n^#��R��+Ah�s���@�y����VU/t��?/�5����|@�zS�;#�+F�~�������~����Q�jdgj��8�)L��v��.��! �<o�E�>����˷��g��#�=�Y��'��4���w$�H���'�j�#V$/p�3���6�*;�i���.�"w��Z�5,��j|n�_�T����8fOs��M�(3�kC���8|�&#?}�6��y�!p��Q�gg�v�tZYg9�$�75�f�Ǌ�����9xZ��	�|�M1�=ɕ?�GZ�������c����B�;u�?Mh{r�g����ˎDi��E�0��TM�B��a��M�&l�hĎ �����H������fK�vj�* �,c�O�j�7arU�k'7�)�\3"Qo���?������D��#,<������-���:�B����9 �.���@�p]��s�b͸�dY�����>��Tz�kbkX"5US�gZci�N���ӭQj�Թ���h�=���7E`�q��p��bPY����oGO��(L��v`�6��䫏�Z��1��~ݔݩY���R��%(R��l�}׬k���uw:ٺX�:�>��2�ءά��=FV�D��W* Vo��y������^�E�N�*2�9�����@Zzvy��c���SF����am����CPVBF�����t"H�4�j�u�vjS�p'�[=���.@��q[�R��9#x�V}%?���/FVY���S~H̬fkE�^��D6M��	���E�:�&{s[ 6��۾�h�3p[�S�]��Z��[�i�ű�g&7���Urh���H���ڂ= ?�����Vg��������"Åm����":��_�����p���	!''K�1׮/@m�-pt�!&n�'�����D��j��k88��x�v��h,\7	��sfr��i��D��˾?H��4��܇xjY��\�iz�W�vE�9ݲ�{J9��H�$�Ak�R�lQ
�SK�o�Z�<뭻o:�6��G52&��0�>�յ��x���dt d� ����j��wo������3�5�[��y���P�Z�'��p Ք���f�;��۹��t�2>D�kE:�B'���L"�|��Il��17�L�O����ƽ�J~��Y36e�[�l�׺|E�g���?�	p�Vf�&F0������J)���D�E��S�#�fǽ�Rh����I��̀\=��0X|�/T�;h��H9��-e���0���@���7��*d	w,��:�>����������-�.����|�w�mʃA�=�;S8I ���K'ND�e�gd=]�x�m��i�[�lx��F�nl^��a"�F����vsbhYþ]�q��a[��VQPN+=�	X�޵���_���)'��vH����7�cΆ�K�>�V�)ey�Č�o�2����MWd܄�"��,zۢ1?W`�5r�_7�Ϊ5������J�)�u�lS�	�;�5�� V�)�kv��C��O�f�]o��)~�;>CU��vڻ��J6��q��S����;��zA���?yڎ�we���Xj�4Q�ڦ&~�ި�90(�h�f�{(��?��]g���5Q�*��U��ʜ??��Jccr�h��aҦ�x��~�gt1��Fg�jz.��'�{ʬ��^�_+W�,�b7���=p�W3��^���$����V>3S5���vr���U�y%��q�����z�2����ǹH7�uN1�Fba���S<b�.J�uMa���߻ ����:u�S�{7Y{���.f���`mʇ������=��A��Њ���J
q��wl�<��+������A�^t�ff<��T�̎���%d�X�܀yW�p�v+�Ƕ£#>��)/��c�*[{�օϡV{���ȴ��
i�O�ET��*��|m;˅OjK��0fcKW�<��n�kl� �'+rT��7t����_�ţrn�� ���0���=��ݟ�!�Xj�b�`�CgY9��"�-|���������~q�����r E����YW �b���z���%��.���9O��7��_��.:�,�7c�ϟL�U�ȅ.C�Ӷ��$��O�%c�7<�Vc�v�%߰��p�L��{&���o	���_ؽ��[��Kك���9�Fا��@��c���e�DstG�{ư�gw��_��{mM���:5*�Y�8�X`�(�Ӯ�����.���@B�>4Ikm��p���g}IEǗW�����x�� �pZ��F�[o��!�`����[�l��C�)�R��A�պ��7?E7��rzn�/�j�=Jv%K��i�O�y�����a�؂V�Ի�ҙ�M�X��%ZJ!ӵ��=!^	M�f��Y[�|�ldξU�<q�gT%��$2��*0��s���˜+T|gB�6�g'�ip1��}ƺ��m���d����W���.�O�j7G�����Z����{���B�\^�rM=��Cc��Ձ���jM����?���K��.,�,��h_�Y\��z�W�8ɺ����� �{�<���4��9�~@�q���URO�0�	ˌ��z������;Š�2��=%Yќ��ձ2�2�΀P��"�$���������5�ދ���G\���1��ǿ����7���f�p�xc�����/o�n���4y��s�5P+�)���6��l�K�����cs��ߡ�Ѝ�6�=�*iS|w���Qj����P��oWk�(a���WKp�)ҳpsW�Vd���aÆ�hq\��`�!�wNʨ�h��U�e[N�����@�S� ��=*o'�� ���b�^B˅ bk��7���,.������U~�L�WT�e��z�+���#��1N�uzB���T��h��n.�z5m�3&^Lw~Wd�!8�U���t��E�@�n�^,�,Q��������իb������J�x�7e���\h{,c�����9�9��P�(���
.���zb$�k� yﶍſ/��Ŋ5�������q��x��ؿx� �/u6� ǚ�b��G���k��d$��1��ץ�k�����K��EOw�N�h1R��{kl���ex����7�I�*-�Z�)6'@[LY����?���r�mj�g�Ǥ��G��i��kE�|�T:���/��%�M�qPH&u��Z6���5]�rS�7nu��]����a�y]���^�C}^�Eعc=V��<9l�Y);�MB�6r���vb���T��&�9E�J�©��j&���t�di\�r����=�J|���E����x�;.���~��z�F��.�o)*J�_dTy.{��!;k�tX���g��o�B,w8Tz8�@H��m�f�DڍN�cbE&e�����i�o
IsM]�U�\��سmҲ�2]&b�.�?�l���Tٷ�+��RXJJ�-E2��]�'�i�����a��k�I)��+R����*�m���U�3���sRKi;��)���O�N
AWG� ��@c��ހm���-�~�cۋ�j�a�MW<��1�"��-,H'���	Ei���±�s]�F�ܟ��y����C��8�&o�N
I��_�M����:�ez����lmF�Z�C)���[)
�Pt�lP���┠Q��Ă9��K�a��1�K�H�������Lpz���:�L��tƽ9t��%��C�߸�C]{!�=Ek"TG:��ZΦ��rcu�f�� �6ᐩ�/:�F]�ڟ*��triih���OD��(V{�@�2���Lm�Ӈ}��A�K���
*X�ol/�e�/S�K7�׭�z���V�ծ�OKA`����Zs��I ��!��Hz!��<�����H�rm}����to�E��=4��e���E�����gL��\�03:A+�L3AD"�2<�}�XW�1⸷�_2�ݪ�&����
w_�P�;�Y���i��F�ˢ�	��7�E����^��r���ګ�ā'���/�eǁ��f8�ڝ����r��.�����Z���=}�����0M	2��yW�+|k��q��xoD~�����6b;#a�����3+��%����xc�b[r��R��M�]�з�NV;a�ٛ�q=\]w�ţ������Y�+fm`����L�|�$�u�#E�ޜ�<6��rl�s�ec�}T*s�4IO���%+�%ݗ�M���*.-|OWgs˔2?:�.1	�T��=���t�Բ?m�g��r���JPL߬�@��$Q��&�D�,��#o��L��~���S�ԕ��A���W�Ç�%��x҆@�8����<Yfd�6v��� GS��;���AepF̔iQަ�}w�hnT�	T�;�k�O��My{5X[B�O�c�o��H��� �o�
0M��^���I��ɟIj�8��IF!��jMUu�p��nc�>%�6��-�t@�L��Z �b�;�:���� �i�e�R�G��A�F�'r�k��a�g͍3h��ݘ�<T[.�J[m(����������
�ݷ.�m�kڅ��ۉ�;K^r�<g/mH	%��Vsk�L?K���ʓe��N���Bဿ����R-`�)�i�W�{`�Q�zS"�a�2�h���/)k2UhxZ�Ra)+���ܨ/����X��'��Z�NmX��Ewp���9�"�o�gy�E�w�5���&�����O�	w'�Z�s^�B���L��t��|�J&�;a+3$vXzh�E]�����fM��u���	[��YJMF�!��"�r��8n�[V�:�S��Iy3�t��nd���{���b�2z�CtP�_��߰�_W!1&!΄�`��3�����e���UHlf˲�������.��fhj��k�\�}�@n^�u4��z����A�I"؂�+�3��ݜl�4�~����u����+hW9�j)fV!�SC�нv]�誔�����%$afh��VR�c'�O����N�"��+����M������p�q��Y��6�ncJڭ_槂�}�9�V�Wo�44h��	�񜉘�J�POCw�7B����lE0�9p�[7�d1��I�����Al3����0���R#���jZ�M�D��zp��
�]R�s�x@Z@�]n|a_/#g��	V��,E\6��qh�ݙ���q4�gN�!���#��,
�T���������V%����*�݇=n2��d�{��0
�y������>
ޟ��R�yV�_]�J�����!Ϝ-�g�Q7�D��8JQ7K�6��q�V��x�!�o��8�FąIڕ���WAV�hx��?�u���\F�mv�$f��F��fZg���ճ�^ת<h[#��#�"��'�:#��l� O�����\^Wl%���"=B�����@e��t��k�a����j����2�v���JŖe.1��:ڹlS���<S�q�ߺ���f3$7b&
��?3��l��V��^ͱt� 9v��H�T'��t��Y/��O|e�)�;���[W�N�U�WoMh̘i��&K ��F��M�)���H(V�~���w+��_[ ��!f����쀾���p�f���YI��Fl�ވ��'�Kc�	ʵ�%i���ր�j��d�u5}�|碳���\@���J��bm��p�1�ɇ�s�ܺ��S�&(*�H�-)���6���"4�T^U���`ɗ�mL�-�'���w,d�5�K7V���|�B���_)\b�c9LĳK�#�%�,����k&x2��PkpqEж��y�u��f�a�Qb�&
�{��v%���/�w���ҷt�/��I��o��������/���'<�z�w�?��2��蝿|�>�?�_U����GU�U�Jw��-?���އF㥮*�����PK   �A�X+���  D�  /   images/5cebb09a-e86f-4cb2-800e-22da09d26481.png�yTSW7k+u Z�	�5�����dK+�т*�"�2$�!L�
���QF��bŀ"�@ ��IH��D÷Ͻqx�����w��ֳl�9g����>7湴��Dz��EA���k�6�������o��*���>?���=�'|^H�{؇@��A��W{j�<\s�W۳6d׳�c�.*��v������E���/�_K l �~�i�����n?=~�d��y�>����g{�.߱�k?����n��������k=.����yAʶ�S?7/ot�Qi�y�u�̿�]1�����_y�͜�~��z;f��ln��	�	��To��*���w�y{YJ��|���\�wr�k�0�g��2)��@�0��P7`2E��]��Su����\�64��b�BU�c�C�qs7E
{�U����|�
d� d��\�դ<M>��ᖼ# ,��m���/;K�5������k*�pnyv����ßM�GV�m�o����߆�6����m��m�����	�(e֚�ܩ�wW�^d�����RX6�,H$}� �o�h��x���X��p͎�Q���cNKCnBI�q�=qHi�e�{O�1=
x�k��U���m�n�$[G��3(��S����(WX�}�O��	��@p�9r_�6���9m|!�X!?��5>B?k��9���<W{���z��˿`��o�_� �ix�2������{�7��k��{����W��r����BE�z���V���7/��e:�I�ېc��2�?�)N�oL	G

�������/�O����"���<�Ot�"�<��,�z瓂]ǿ�ϡ.K��l�V)�8K>/��i|bH�	��w���*���w\ &�[��F��Ld��4�2��f@O���Ӛ�h^�d�+��K�������	(��S�|M��;) ������F�gAB2/	?��{��8y��v�BX�-���"]CY�����i{�\���D�=��j0���f�/q��!������M�u��>��)I�d��dK�nɁ_����Xދ�9s-0`�R�c8�@@�5����5�/$P�]�ر� �tZ�J�+R*9��|@\��5��v?��>���:��:���$2����Lb�z\G9��~\��.'�ny��!��-�q1Ș|B���_]$���	������|oS X&p�mW�c��~�?���{@�9�(���uX�MH�-�0P
����`����$/�������1��1F ����7r)D�v�s��Z|;�\h�D,1W8���gƚ���8f|��J���W���~!Řn�ŵu<��K|���ޔN�]�.�v-��r��7mrue�'q��L)R��+��¥�����z��ϑ�g҄DM�f*�r�Trܒ"S�+�#�+����ϝ��f!(7@?���9�#�?�}�+�a��כ�+��EL��\��&�I��}����I��]��g\B��Xe������)=PI�Bc��<�p��Kb�DB|~_��[$� �Q��=��g�����I2�uC����,�=0�����霫�3h�����tG��n��!�Y�^�&��~��"}d�}vxf�=<���:�G� 1��3���`�}n�ϴu+/?_��nF�޵��D��x9��k��K�n�i��+�0qa��1�y�8��h5Wb�م$59��C4����.��9��ӀT'ɛ�<�T�/�'6����~�򼚄��)�YT�\�	���)���/(�Ye�� ~��J]��*����-M��3H1�nlش-�{	0�`{7i�$�d陼'��K��R����ԣ�����]�QG��P.N���2��;��/��~%�mRN?f��
���<�WE�s-t 
��v�Q�`��m���4@FfUyrv?�m�))������-�����2.nxJ�Ǟ��߀^OJ���X4F�M 
�m%	maz��k�j���O��� l��fI_6.;�G)E=ΫM���/N���쳰,F�Z �z؅�n��?؁��< ��S���¤�h��Ge l4������,�nY)����i���8���>c�7����x&|Ό~LNߖU\��*��9.�S��(�5����^����@�Wǯ�*�Pq��R��ySL
����oâ�z�T@�� �ǯk�.�)�kD�G�e4o�����o���UT%+?5�DO�/�pƁ4����}��"�sS�b,�B5�/X�ٛ@Gr��!y�6��ē�M8�7�I U��� ��[Z��B+j��t�|�2s��R��I����;v���Eʢ:d��ЙT��ob���l�}/!�0�_P�u�[��gߊ2Fu�܂Y��.�T�����f�>�g�?�nY�������g��Q���D��R}=ax(�^~��?06����G/�v����p}�37���o�����s�"e��X�����z�l��cZ/�)<�u,D�Sܮ�E$ �CWL��U{��� DC/@���PcA3��$Z��{7�(����a�]*'��� ��̛FP	�g�G��S]D#=�
}V��.=�칵oL�\gɤ��Ìl2ܚ��N���i��6@KI��7U�>W��ʷ=�i]����Y�ݓM��[�{���ީ˕�ח�>H�=/@��kg��4�|*πTYU/n2
9��֕��^H����.̥OL��&�I���{����]��Ш��k�y[���X���d*���D؆-.*��}�l�U� ���Q����l�e��e,?��b]D~^60V��4���Ӏa�̟�SB���py1�OT�78���-ߎ�5����Dx~ء�,>@�jeSҼ���������rt*�s�!�[ͧΊ/S�F��x2�A�G9P�GT�� ˞��@���'��F�L�W1�u�p�X��YAR[,��8'�$ 2����0��o�=�
		Z�/�dvWC�O���{���.Y�4w<Yw� �Ke[�v����˝���Y�Lw��^��5oW[����e� 5����a���r�/��Rq/��.!�kV�����#��W7�h����S��k�|�Ю���)V����<+KbP��i�,2t�=7�����,g�r�S�4�՝j؝�&���X{L��^�͝�H�����浺K��,=t����O=��`=�k�i3A��xM�t�y��W��^�����O�gﱦ&��~M�pG�3a��f@3H��qo�[΁���ﾡOm%�Z���53�9o�,E�aXĿ/����Bx�_f��;>�B6����M-'�x(���];��k6*3�y��"�ץպ^��r��r8e:��M��%��G�F��E�Yӯ&گ����/�Uk�_祻����}I��hi���2o��6�^��_7U0���p�<��%�?LD����л����g(������ ~O�./o?r�}��y�3��Z:V	B6��U��3A�u��ʨd�jD���\�Κ����ӓGv��n$�[�l�} Ȉ��H�H�m�O[ó�3MI�n�Y~X�������F�A�	5�h*���U�k*�B+�7�Ŕ�(����YY�ɩL8d*Æ9ߦ}Z0A�O���N�'���r���Y9S��wnC+q�������2�>��N��R�5y{!wK��(��x�Ӏut6�^�d�_&őo;S�M�wQ���}傘ۗ�v��?�����=�2�ϛ�J2A<�#��nV�x�[��� ���]�9�]��z���,�:���Llʖ;��� T��3&�_����^T����2ET��q��N����9}�O$�[��v� �͕�,Q�̶?��܂�Qp.��8��uE�B�%5�X��nb�W��j���MY�"���U?~ j'�rA����p��&�7��,�0�Χ�K�P��sE~�*�ơ��r����ͬ�?�Q�i7��̏��:8�H�2�9/l�(H<����^��#�$;�G�z\���,��t��իޗTV5���^���l���|ϝ1����v3�[�9+�je�ŕAc��hk��R�����'@�h���FM��m�	[�b��`��baW�a=�((��2�or'�T�9�pZ����]X��,+.ˍs@+�{e
V�K�n�J�5(�0��P�$K�Գ4z�����wK��nO,!,�N����k��SE�j_��ƞ����z20�kT�l�3������}�{���R�A/=&n�b}�k���8����f��YŎ��DU�?��n�����䐻~ؘR� �j�[e4�;:�ye$"�C�w(R�3�o��9���{���=��:�6"��x��
k3������Ṗ�ɑ#p���ͫ���?12�^m���'t��2A�f1��Rf�M��h�	�D�:[�����h�:���p��>E�JuY�p�*Cʇ��;�`JLz�4�e:2������˗Fb<�f��+��J�W�UG%'����j�����Âq�l�_�τt��@ς4�A�5��|߄�v����61��Ϲ+7�[�,���Ώ.�����}5XA�)�X���ޖ��4TMWу��d�2?3.� j�!�9���~+n���rM�MG�#Z$/�¢	cd��6�}�d	��ȟSd:1��l3fN� �d*O�B�f�sC��g��<�}�=�����^��Ct���]�'��$d'�IcZ�3�ӧ鑓��nر��؊@*��i�5YyrJ.]�2$��1?��WJ6��C�xoz�qxO��-^�˭^>���U��d2�!��ݿ��5�i�իF�'��:�fBWE�撈����s#6s��:!�Xh���R�!4o����I�g��5���޾oW��"�����(>��F��=,O&��
�ݱ9��4(�t6���8��kO��}��l�뚖���B�T�@�I�|�>}d*�HUd9*�9�p�ԂE����7�^>�z�u��m7�7��;8��ksD��%����B�Cy�90�0ϲd<ռ�X��A�3�v>{��1�aEw$=�%&�S�o�:mW�b�:zs�LNc��j+����c��e��O@H�Xi�8��c� �W�$g�9�#����1÷o��&r�A�.��j��=g��MV�tSjy����ѼC�F�/�b�Q�W�@��Gy�"�Vrzώ��Y���*�6]#V�a�G���nP�^熯fl�(ǻ %��!`K�����"�{jd�Zw�8��xr�����
,����?�ԓho�F�rwc�4�c��Lb+��F�P0�[��2�P������M�����>z��|�N)OJ�eM����7�E!v�6�S�̕�#�;�/�q��쌺��}��Y�v,p�W�d�R��F��x�_�V8+Qm�WD��>X�*�wI��R��\ϭ�}𺎌c�Mu��2��c���n�L�;�������HQ�Ik�mS������ғ��*O������:���d�oE� �OǷ��'?�gd2��[�^���3�*i��lk�G���F�҃S�\�G�L��&�ۻ��u) v��h��f��+�T�����o�"F�_�ʤO�	AP�v����<�9:�wk���K�=�X���@�ުN��{��`X+JP5���ϳ���F�9?�U��a�4�R��m���f2P��Aek�0]�"z?�8��044����t��s���93�}��'bz��!NB��[e�zN���X��7"߂NaY�I*�Vj�c��i38������0�ct*���4��s�J��a�ݮsq��'��}�3���vO����C�BJH�LIP1�*OO��ARt�oc�յg&��X�EO��}����%C��dD�Xi�ዪI�|�lK�ڷg�sĺW�1���S,�xk ,X���,c�ޥŦ�c��K��=����a�}���4Y�v���T��2>��7�KX�iD�
NV��ED��02S#u=�*���Ao5���� :9�/t�����u������}K/��5��y���U�L�mt�>�K�5��'ℸ�N4'3uYc�d�г��H�rAv����9G�0�
y6�he���:��l�Z���?l�\��1�R�a'õ�(�������-WD8��̅�8p�s����dQ��-���G(����5o�����Qf��]n�"��p�7q��:g�H���?YK4i���]�4dQ�ץ��U1<��;�G@�d�x�_�6_M���'�V���r�e�����_���#_,�i���5�N��YGWR��?�O�ׁIVeW�9F�s�<mo�#\���&e��p�W�^���ź8�5��כ���CR+$���k��y��nWx�p��S�i�����7n���A�g�X�{���g��5j�����C��	")x���H$���[+%됐M����i]�%�q�j�>iꭠsނ�<��HV��OY�f�#$d,H�} On���Y��� ;g����U�ae�,�A�"�I��՝���"��ꉋD^�6�;�_zeF*��r� ���P�9�{��� L�F�$�h	�G�N/VH������%��I�^A� ь3>%9���^�;��&D(O^Ȓ�����x�,%iis�������?�elb�5Z`�]]u�[�k�N4�YwR�I�k6�Yp�C�%����$"i�u�����G��?��ҷ[lւW|���. ����Y)G�6�w�/��>�b��5�1�k��IY�#�svA3��~3��5�'�3@�_�e��!�G����iI/�d�O�
�w���j5�	�~�����'B��:�g�gB�;�u+��+Wʽ����T��%����ol�q{!~n�E=Jv���(��۽tٗk�:Bo�^�~o�*"�mL�W ���l������z�0_��ܻC�̛!z�sn��iV�C$3�Q��!f�+ -�ˁ[�d�Y���|�FS����7�����Ր�>��vv[(�l��A)ØL*�]�������&��xRnC�"]N8�N#F/�;���d�,x�B��M��Mi����M5w���(�p����ղnR�뒧U�+yD���::|,Zv.�h�ic6ȱ��v/�(��z]7�����F�F�}N�U����A=ą�Xaӝ�J6������=d\�����-��W���x�]�A.�-�1��p��Fr��-n�0Hb�Ͻ���e=��XԀ�|+&+ł{84�<�6�Q>�#`�m�3g��l���G!�Q�U?�e]o��{���@��a�+�e�p�)	�L��ҋb�1c���0�<�'���=�I��뾥����;����^��U�ǖ@��U��О�,'q���k��t�J� � 6���r�v��6 �O�&�+lm� �lTvqb.�s���|�<�����"+�Y'���>�W\�o@��0Cu�[�d1����<������q0b�����-��?��Ϗ�E���
�W_���ui��(܅��"��]�n��
��Ћ(&�/5U}� ���?��Z�?��̙.jP7J�}3�x�ţ�طKlA��m6�9ѼK��d+��6l:k/��hE67ѝ�����QY+��6ő�_��MK��_e�_��Q���j,����+i��<"@>���P��R�t?<wφ��L|UkV�	Q�Fу$^# w沼]���CJ]�Qy�U�U�	�Tͱ�>f�=���J_���~�e�m����Q(��Л��å*#d�)�e��8q�7��[lϕV����b\���%�s �"���/�:L���B�ܣǏߓ��:xj��>��_�?���Ri2�W�&�|�֖<\H)0FGy*#p;�xq��TE?fj��$"�����#
L��|�et��4�
E�zص�f���;k�ʦ��yy@�a�����"��X��y6���	�,:9������̼��h^|83C*���'
Qc�˝ԃ<�S��W�Tp�d89JL���#sޯ�C��Y�G�_���C�Å{'���!g���Wa>PӒ[!7�Τk[�s��	Ǆ31ѣ�%� r�4"֖�%P}3�4wo�@!OzSn�t�?jۦ"��!`�U;�Hٺ,�r3'���y��6���k*�Ȑ����� �N�����o��*?��V�K����&���"2�>=2������x�ꂝ�:�'����T:Q���{�i�s���;!*�ź���2;;a�E�>8���tV(y���S�#�v�N-�Z�:�7O� ���E��I,�ԆUN>5��n�U�١��F�w�����s��Q�����'|�r��l 9\�=�]y�5�c=�YsK$�N��0��݋���ħkn���B"y�77W��ߘF��2
�,i�5ֆ�*���Z�*�<߄��0}�Rcc<=S��M_�c�y��U$�e��v�}�����4,�ϻ�ɒ�pB��c�u��+ƶcw�̀]oKQ��ȱOUQ��d�Б�/�5O�N��O�.V��ѯ���簯28�Ra�Lb��ֽ���W�d�*#2��+{�+h��u��g�!y#��;����h�#�Q̖4<׌
F.z-we�>�]D�)j[,2a�0S,�����"�8��������)t�;����8�	�J�ؤ'�{���84��{��4�X�:u}����@�7�`U�2[�7F/��/��,|�M缀�F"uK���x�Q���� @0�Ǭ���2K9��Tj*���V�{R�!�X���Y��{Fr�}������҂9��z����*m��'V�u&O���07C��`n3|Q�JOQI��L%�᧥t�~�H*`��Ah��~'�߃`0���Eu�Ƨ1��v��B�y�l� ���v������Ij��&���:��V �AV�D�P�Kb�2��z�"9$�����#�l����T����EZt��n�:�O�0h�W���\}!�W��*�mXA��@r�0������߻���,B߳��G��P��\�U��_���ܝQ�p���Q(�LuF�1];��'��WEK��M�u��� �o�Zՠ`��=tt�&-�o��w�k�b>��ԜPQ"�V��N����gY{��֧ؔ
ȧ�ﭜ��%�y�5�LNe޻Lbx�M����V��qs�������Ѯ�۫,�Xюcok�$/�����'s��3T�R��Nx��Z��<2w��һe4��G�᨜����JWE�z&o���ס������<u�-g~�S�w�D	�����'	(�Mb�2np8�x�v��@|fO��NM8�'�9�Ei����u�f�\u.���u����M�c0L��3���\�\��aw*��~&5�`��`&�X}Q�@��)�ܰ=�J�m�b/�-?�f$Ɇ�є�SYVg��5�V�Ƨ����	�����T��W���ط��9�^K��\����7q�L��TqWS�0�9��]��6��~f���/���t�"":��.I"�dl�[�J$��pd����q�b;��[O���&Z<׭���&���\�L<�\�>@ՓG��O�mﮬ,��7���Ń�r��L�mFb�X��n�+�L}:�e5��7]�]k��u��;��������78��M��A��(�~0������M\��׎WaZ��?�k�C����%�S�������j�\� �e.�A�ͷ�KN�^_�?�0�l,ۊ���?4l��;��s�������c�!ǖ>������W���46�d%%���6F�M�?�=�&��GJ��{�%���m� oY�+u��%�2���ލB���O��1/�,B~�8>V�ܡ�kVZ����y�I�jnk����!�Wu���Ti�l��nz��Z��UUAe|���T�iw1�����ޞ�&��G���@�W0OltUb^Pc�0�;̺���:#kC���ix�f@��&�um��1H��������$� `�&'CrP����	����4QPn��14;�1�<��w�;'�e�=�`��y-�����-�o7#� �\�r�i��b�� I��b����eD�W5��;9�s�����EF�GM�� ����#� �苩F���w�\%�����.�5	y-����l��i�B�(�YQ�� ;�c�����l�bu�ȿݾ��Ǯ���t׼W�s[o�m�J
���G�6��Z*���EZ�BάS�%%	N("�}gN���iCEW����J�O�c6��iK ��E-�����|�P?�H�%�$_ѺoH�w!w_�R5�!s�'��M�:�&��`�D���VG8�$��{ �'����B���W�.m��x��&�T�3�I��)�ÊHg�;>X��/�M�
��7���Wj�[����AE���`}�${���DG �����]��j,E"�����}:�R��ԡM8��w;X#������]�g�Jb%�:dٺ	E��� �V�e-������M����z�����WM"zl0�$����V(�~��!S-f"e]�q��Asl �}R'łO08ZJ1ʣ
���^�h�����!�*���#�s�-��R�o�껡O��1��BS`��i�Z7\W�,�h�(z;Y�/(B�V����D����~��O��^�C����Jt��H��`��^�UZ�����A�vrHE��:��*�Zl��=F��] ��r97
�{(��80�U����׬���2+UQ�,(�dGlpn��Q�^k��V����7�)���B��Ƭ}��0�I��L_qBṄӃ0�!]���Q��<��)c4J�\D�ښY��
�]��{��&P~vR?�u�hf�/gw�>��6��e��i,y����O$�����?�6��Hx���7�۵�ՇYf�(;�Ʊkrb	��3І=��Ё���
�1�f�s�N�+y9nͬ=��jTTEh9gNs�:��Y�>��n /�rQ�`��ͺ�86Q�m�O��F(��,�abS֑��W����Z�2;�@�M��B�oL��WP�s���HkH��Ԙ/��]�;�)F��DA��w���ς4�R����>J���8I%vU�\��tY^���������T6=:@�貊<��ޤoD
�Q梲����=��\������Xw�n��yb��{��[S��X	��<Z.�-Uk
��h!�4Zχ3y�Fo��q�㎠G�[3�#���+m����r��g���5)��eu[���׍�O�{��˄��ǭk�H$N����=�h���SA�p���x,,���'�;�S��o�mIɕ8� ����^��I"*�
~�#��`�7�K(���Y�*AD���sީ:����B�Z0�K����~w�~w�� Ф2��{g;N���i>�g`Mm��d�~�������W�޹K��2n�Qb3<����687��v!�Ȋ�nǤ��(����@�W`ʸ6���ŕjl3��U�����W���q�*(+z�C���^�I)1��iQ�,��9S�����7����?�6�iJ�L&���l.���J ��IjB]��Õ��,�0q�4�ĭ�3�.-��������ae
DX���$�-ޔ����^��&���Bsu?�Wʦ˂�a�ll��Z��vL�i����}��J|,���?,;UA��DW���^%E/���/ l [Z(��h~d�=7��1�zN;%���u^KR����>�;d&�S�UVi-���xlJBW��S.�1��NUR�s��9�'Z�C�F���$��O��M�$��V!�jeEH��9��VHܲ�%E���[2�nR�ʈ�w��	@4b�����a�>�n�hY1�$y[�>�����V��$�!�$QBv�2�2A�rkT	�!	��Zx�v��W��W�f٤{O��l�,��������M{�X��z��T=������f,�}��Vc�/]Tb���	"��O6.���nv�4v�93��m�H����O;�7(MBR�u��?2҆+�w9��`���x��T����z���n�bk��m���}����v��`�}km�+�HP��ڵ��mbW,�ųQK����VΤdطC�~�1�й�z�u��2��#u|p��c�E
�L�9@磝_m��!2씵�s�7ǒŋWA���n�qw#��,x?����t�N�}�TF�pi������A��U��ʳ�74s��g��o�	R�D��R��]+
�3�}v�vG�.�KRTl���D�:77{��)�w�<~��j]Z.Ҋݚ0�t���^�^�"zd����	�������k��F0UdY1Ɇ~�>���p�|�b���R�goRv�R��R�h^$˗2��6�ȳ��RQ�س2�L�0�_��l�*��|tW��E#�S�ÞX�:����#�!ǆF��Vwl��&��[��uqd�x��kU�Rk�m��1�W`�ˊ��eww�E${`&隧/��	+zm��${Qa��A��qTζ�߿��Д9��*9����'gH�_��@���>����"Tb��E �U��܇�J������#M���D�3f�3$�y):�O�qh"F�lo�5�(�� �{wD�PK;q��7fN�@{���h��첏ަx�TO�&�So�;��_�����[�L&aP_ҰP$���{��p�E�fr<Eg�x�VT���]l��D�����V�z4;��pi�bѲO������dβ^�w��{�hrm�(e˧^�ٻ�r���B�7S�~Is�I�fό����{oH�ʵ0[���?4(y Z�b~��m].ت*�"|�����C74]��Sf�ZB��Ѡ��j���w�7Hϑ�`	���=�7���e�
*-�H�l�l�P��}|��|��ݽ�c4w���]�e�e��3V	�S�d��������������U�gz�w�o����S�ߕ�C"��?m_~�F(3FlF�9��{��Bf#��� 7�_D]]�km�/N� ��G�����5Kn$�M??X��,m�h���ǆ�#LQ�T"��$2u%��W��E�¼3;��%���O�>�}�]��Q��k��rU�w�~�ݿԠ#�Cm�&�΀�gb�B�N�ޤ;�����
����+9��)�T]:��pt?	E�q؈?]l؋?�!��y�/ߛ0TT�c/���^9
�����R�5�n�ry1Mcǩr�z~,>��u�(7@���.���>>�.�>dﻁ�s�A��ό������;GN7�I���x���(����f�0|�Z����6��tP�d+�9��޼��`1"���_t�[���	N��-�a�ￗ�?*��i!At7< �_���C��"#����6�(��Ձa�o��,K�#�b�_� �s�P���&^ V���� J�R�8�?.��n_�D�
D���h[����{�W���[���h�J�*��Կ��9x��P>��-\��rMΨg�,�~�g�$^YG�@���4d�(�g:�@��O2���8S� ߳���ë��9]�L�=��C�Ps�>%#���w�h�VV�$��p���ҏ���ύ�����[:E�g�A��qf�f���}���ݧB��� b�@t��;2�b����m�'���e��Vf����C/e�S<���B�p��`����'�ϋT]����i�y���+J��X=�:1�������6LG�?+��ڗ7���p�QL=�|�-�6~�Sa�}����?h��qh,[���T�S�QW���Pg��|~�'�ʣ�J�������q�M�I�c����L/�]y��������ǣ�K�ZxIk���'/�����'�g������ߔX_��&Z�Mkwu�i9�;s�JMG�K��3�{}&�EcZ�˃��	󗲏��v=Z?X3���x�7�o	B~����d����fvK�o�*���n[��R����29�4����df6�hl���r�14����	����'�(�L�sm��:�&�l��it������k����v�W.�|�,1:@�y󻚊�[hY/ð:}�k�m�ua�r�ע�\Ӽ�O,]xb>KM�͸ߘ>�qg��4��aW�;S��nq����ܾ��6��D�H�Tu��F�*�_��sA|��N�o�.��.�!!��;��LrI��� ���q�B��ɺ ���<u�D��<ǘ����"_
~`�>�'"H˭c�e�$G�W�0)�Ȭ�������<Öz�u�����Cu3мΰ1�Ÿn��5���笍���Ź�h���w�\s<�v��C���_(�]1!3�U����nv���=~�����b,EU�
�cDg�
cIP��"���<�Z�Yu����½JN*7���|�$�Pr��1N�����\, ���^������4X�ZO[k\7~����cT��|��{n"4�v�I�'�'�����ĉpn0e��y���XP����x>��Q���qi�/Ђ����d�Uv��k!�_I�kj�?���)xH7_¹S\ëU��`��\�p����#/�Eg��n1X��3�e�ck��ԉ��f�gic6��.ٟ2݉�����]����7�(k+���S�l�fΐ��f���s�N����	gh.�c��޸h/�B��v�s��WBw|ǾU���Sx�h,%j�^��~g��Ժ�`ڃaRlͅ2��;D}p��������ɡ���>��.�,F�v�)�K�i�b�%|��Q�2e�f��	�z���1�������r�DO�@��.Ɲ�Q�/����⿭	��}x��nni���lY�*N�	����]4�pt.e��3�/!���(V/��n:�R��X����1�K�����#����B,G��d�`MP����4CO�E��C�
����J�6D��&�{7�������pc���4v�(%���+�Ldx
��^	f��,V&�^�{ɸ����ע+'8.�f�ܤ;K �~�Wf�}�W�g/4�;KQ���[�RH� o����<�>��c��H���u����o�d߳C������N]A�P3#�D���'�A찌�������W����]����Pa=_hh4nf���I�`�Zh�ë�+������nC�>+�н�?U��C���N"c��JpZ�5u0�Ĉ�(�1���+�*Wxx�g�׽�A�Y�Ln���K��K�N�i����`��^rd,V��[%��ĕ	�串>��p���)8>5��~-��`�[��_(R!�!Y�G�j��.�
�������&lдzq�P�������H&�zЕ�l*��o�V���B�W��@����W? i�D�ME�A���*���9����T��U���u�ش<�B�	��'��hT���tV��%m�0w� U�� n�	�²��:lΰ6��}�>��Jc��P-�趁ƓPQ��j��24;<�쿁����Y�uN� �6�n2L|��c�Ze�������OyJ�I���u"�c�N�aϸ��W���
�,�(�Qe��9�_=�7�����X�	9��������r��w��o���R����)�ܥ@x�z���J̐uxn���>�&�«��_���Q���)�T_'�����,d��sDK>����zv�ܛ�n��s�!ӱ���V�Pgr�����b���\1u���*������E)�A������ȹ�öZ�v�
�wc~�����x�jpY����G��]Y��5ٓ���=�dӒ��#A�_�gWʻ����p�\�=�~��[�B��xZ_#��\;�局T� 𭀓�mr����;��"w3Ȇ�&����G�{�Κ��vS6�=��!�D4�uY��8ס�/8
�Bk�ˀ�"i�C�e}��M1z73A|Mf��ҰY�z�@y��nc��~�¶� �ڟe�o��<s�|Cs*����r���"�۷^tS����3����&
��P�p��DHA�yj�'��W�َ�/��
R#S�F�t��b�MP�L�Ȭ����?�ݑM�%�>��B�-�����~�:��Y��CFݺ�'�FH��m/���&]�cK w�4L�������c ��:��� ����ox��� �c�l!#�}��χ{�<5YPk���
�&tU�������.*�O��*���0�����G2M��IPd���H��@g
�BJ�'V������d.��o$��=�V�H�{��9��--~���5��p�s<��OA��	�%=7�T����T�Q�v}v̄`"����i����.z�����UiJ�w��(«���q��� �a��]�*#+�Q-��Q���uZ��� m{�ؐ߉qة�i�������:(�*x�j�b�|&��;�_b �����豙9�R�����qx�a;a�추}����s=�{����x���4>��&�G�I����(t���v��$���?�J<A{춤�7��7��YH{��.HQ��y���O��_��قt�������6��%D���1��'E�	���]�
S���܃߹��?�Ci>4W�Cw���rg^��xڣ�v3P�*��LD3����������{>S�Z�ڙnX]��xb��s��Q�V�R	���a)�-�[y\����B��뒔�^��i�ِ=H��PX�
֣���/�|y�L0��#�h�ɁkWf��<�Fח(��SRj%�|�yø6��w���hc��=7����Z�Z��/���.|����Ԃp�-mݝ���:0=I (��D���5�Ѝ���#�Z&~x��_��)��`p`��&(Niݧ����w4��ܲ�o=��9�����TBͧ��o��_�� �Ss>�Z)&�+�Q��f@��VN|��i�a�D���w�A�~*�-%���f�q��] �㷂�uSw��2�ED�+���Rv4#���y�VD����s �`wu��Ai��ϱ�x�8^Tkx�B��&�=rө6Y�hH�P�F�YG�U�$�Z)����ۍ�.��gO����.��ʼϠ�5�7�͖2R�����k����n����?���T��=��h[]@�ր<68<5�y0���H}�a�ƿ6ȱf�����z���_����y�\c� ��:(�2r���/$�Vx0#���Y��ꚴȹ��� �:��q��\%,�|*%��.�_�S"5�����1�K�f����� ab�z�U�w|*�� �G8�u>+�?G�]�Х6H�)��/$H��hOp��tZT��Xj��Q�OQ�rȭ����z�~ss�|E&YF�m��}�R@)�3`�+��F��C���@�A���x�J������o��؉q��5��U�.A�,���O�8�����kL����u��tR�f�C�9�K����Y5Q��f��L�kf��%��,HF���'j?��(�+����JI{�����A^̪�:����>��'�E���Բ�SÉK�s������0���H�6ۏ7�/����=�~W*{�>�B�;z*�?5��zq�v���$UR����BZ�d*�S�(�E;���=�OL�`^�ߧ'%��A|[�V��‶��O�/��������>>h|�s�]3w�i�o�\9:m�&y*g�TПL��ܠа�4�M�v��&��lt�;��XP��f�a�j������t���X�r|$_�XR�3��y�A	~�k��I�˚��g�g0}���ᆪ>�ϝf��#��h���1�4�[9��.�,���c.q=�cQiD�"�:pݹ�Sr��u�6�3���n pD��DE��8)6rt����'�p5N���ظWt��ҹw�?A�6��ā=-�#��V[�>1Y��q�󠎼�Â����B�u����v�-�3��
I�r�Ӯ��[��*��F��#���@�~�x�P��R�/T�d�����10�=?�� �R�ٓ����I96.-271qH�.�vJ`·v&?��{�s2�����ʘ;XW��JR
���L�Qv1�>~8�B��\�9Z�38�Q 662��6����(.�c�\�|wV��y-��1n��8���G�e*��}b E�u}�������eϞ(�L�Cς�&�!��V�Д�tg�n���lĳ���,�EJ�YJ��v��J.���v�ƒzD�����P�q��<�w�|I$28gBf�o m�[���פ]f�P��l��ar�n�ׯ��-���ySnG������M�y5Z�xGZ]-�dP
<s��a��B������tZ�ݙ�w��x;�G��T;�R�`�dW�˧�ܮU�O�8T��i6���ߕ�)R���E��(ʺ�&�>����o�
��A̭�X%� �uϩ�<�)�Y���a��U��L
��a�:l7Q��Ɂ�y0���T�n�0E�����\����t#������k܏7��k'��K�j.ж����?�Q��E,�B}H����&���� 7!�C���ă���]��Etg���7;�)d�ڠ�"�K~I����E	���.C�l��,��@���;�����&����K�8�]Μ39�� ���~T��?��mOj*��hYMڴ��Z����(5���ff�i���7�߱���F���e�ܷ�;>1�����\5c+�_���l��eh�4-^�O�#��R;��MM��,��8_�HߺN���!`���8j��T��N�$��� ���WAk�Y�5�H4�M�u��Ű���������Kdlԁ��R���|-i��p	����4�x�q���O+��s��Ccq�،z8��T��h��3FpP��l-Rk`bbҎ_�VϢ9���~�ف*j�h]@��i�M�����j}3i��.�L�⍸ۆʒ��g���?R����
5�F��SŴS��G��&s�%�؍��[=jHڅׂ�f�%��`��:�V�(V�"8T�s�MA#l"�X谵f�hE�W�q��*`P3Y�:vtkr����x���RvxL��������Me[�����+�s�+2
�� ""J1b(�0#�:��A��Z0�6�U�Q�9�HW1 "E�^"�`��[B@HI�PB�w�s�}�?��|���|��>k���w���0�E ��b�>���f�}�J׌Ω혢H�����"�(�=;)�B�OG��h���[�ƾLÕ�[�i�e�6��!Ơ��LX'R�����L��*���#[ ���(i�@�M�Ǔ�lI����w����*It�2���_,�_qi�������w��_˪�峁˼(�+G|4G���>�5ޠ�Z�k�뎩��ʾA�6�IO��K� ���i�چh�S#1IJG��$�3����x��;�3�f�~�;�H��o�鿁3Lr����a;'�Ľ��X/tLU�:����N���+��A<����N��j�Hc"?jo��\[d	��mp��F12<0�67q"�b�%�)y���|�&���
l�ܨ=�լAY�B��M���M�Lg�OR�tZBC�5�W_��~B<�;�ݝ���oz�����z����K��i�m`��k��ȇhّ����� �a^h§��U��g��g{����7��������vz�ޚ'|��� a"�g���`����SV�L4�Z�b;��]�m�c	(T��г��l&L͛Z��V��݃ڪ��Y���zk}��+-��L�Qj�`��Us�����=4i*�ܴk�L�U�;��HC�Q�x�4Ӹ�O�<��w��ʑ%hr���HΛM̮�>% �䛚����Ԫ��	k�k#�3Ea���O��{q�~;�Q�0�-�J/V#{u�����K�}:�+�%vh���L_e����f���;n�(�3�f�F��W�����������Zx�BWؕ���f�of�q���Ӓ�I�v/n��[%՜/�ܨU4x���R���2�gO�.�G�R�p�ގ�q��)�6 �kY����$٣��#�/b˴_�k���c�������_����HTF��F�<cN�i	��e��� &r1�Cqdۼ�5n���J���7��ՠv�k]+4�_�q�ablxX"��Z�Y�m��uL�&1y��^�r<��Uk<NtZX@��e7������ͨ`�V'����˦ui'�xy}c�s.D�#.�@��U/�g��h�$c+ҋH wt;�2�n��U6� ����|���z���楳"i���3_U�a��ZV��\�Ò��K� ����v7jxdg����L��5�@�F��U�p/Y����ƍ�S�x�4���y�7�1�}�;�7�c�t��o�ε&Id��vSb����;�ƀy����x����ܐ��dgb�a����2Ȋ�[3%��W�v*�x��-�(����o'oC�ܷf��M��N���!�ԥ�YX��")��f�w�:�e���r�pc5�#�a��������u��8R^0lQ��ޮ����>8)H5T)G7m�
5�o����3y�aQk3c���#��&�gw5*�3a��S�޾���Uʈ�a��S6;�[��ns�@U�Bgc�����EbXf�� ���jO��[|%ju{Be�W >P��p�V�G�[;/s����*)]o�>������aL[y�
����{���4�s$AK����c���g*���Ab����TI3�$���$v���.���x�Ǉq����j�"�X�&;�Z���1��=�`7}k���p�P%�=<�ȕ�{�Rn4��|L�$���gMX���h�`(P?����-���G2�{iG��R�?���/��쎥���4�z�_��~(a�%%xCh�`MIG�,�7���B��.�"^s��h�w/�[��4�e�~s�Ɩ"�>�5p���7����kヮ];A�IF��!�`��3�񺒭dT�F'Y�2>����SV��Ǐ�ێ�t+�R#�k˛ƍI�����7�xc5*(���|����ONĊ2%��%��ȿ���K�c���e�SY���rT���\�U������V����"�[_�FӱZKY�g:qhs�+P8�G�
����Qb0�5dP���2�C��Q�z����&���|�ٶ�~s��iw-Xd.���Cp�B��k�y��Wg�z����A����T��3��+F0<��E���3�=�=�"U���� �(6����d��g�>5E���t\� m���;2v���"@* ���I�1��4�	��U�?�Y�˨�G�����*@���a��%*�O!��v�U(`I� і7kh���v�T:�ٖ�g�u|k���l�\,�3c&��x[Hh+_Ur��|������������H�L?#�3�5����mc=
�o�!{���Y3�/*�GN�l���	.��=|aKC�5O�kd#]~��6h������NjD ,-F[}ܪ=*�V�I�A�Y~�]�ۡ��6Ho�@)ϊJ�e#ms����w��є�̖�ϽiM~u_�7�Q�f�C�s
Bd�G�J��̳�1 g�q�wO��湠���_}��6�\�ffY����ؾ��h�/�Xgě����E��,]ZPp�-�@�� BmF>�%c$�j����ѵ_h��dC( �}���v�(g<]��K@<HZC�]뫵uTmP��NI0#V��D�5����7�ۊLTȝ[$��ɜǀ��
iO��%�^� ��oղ�0������.��h�%�'�g�Ɗ� i���~�Y�!�k���7;��� 
 ����Av�c��
�8���N��ϺcE:���ϻ���1ό[I�K���:#i,����My��p�v���2T�Yß��o)1	A��aF�������x<�q��(kU�7D�V	� �M��:��D�^w#�0(r���O�,���j@�
��0+�����
 |��i���p��f�-�E��J��Mɍ��K0j���C��~f<csb~,��xDŤw��1%gp����gd��c���y��]P�2tg|��b���ț�� Y�S��8�<i��M�(��]��x���.� �ŌO\�w:��AO�� �?���h�2�c��w�wu�H�W��3�Tέ��{�] n���rݿ�a	�O��*�~i����|9�>B�#�La�z>>Hr�!�q�oܛj	4|�|����sv�d���#�������J�@́�����;ekm��2@Bu<FK��.إs!��E3����@~3v�~��A%�0@�G��#n�(4�k1H�*�W�Q'@G�yP,&�ghj��3 �W'y,���2����Qa�MĻ^�ѕ�d�F�����2��a0H���#�Z���}w��Q�ڋ�i���e��n����p��砀R[twl�O�xf�մ151������/����e���6��d��,��T�>,Z����{A�}�?o7L4�S����� ��u���Vgu�����z)񹒳#�
��$��Ǩ�mFM��ۨT3��1��o���r*B`�ǩ��l�9� ��!O����b[=�\;�(&v2݉^)�-</�"�e1�E\(��}����S�&O���E��)�\��m�B�  ac�u�bC����7`��Lb�)\�=#ǣ��81\W������� 3:f�Z^9�cw�[���� ������6,'8��+-��r��
��pQ>**�����
7��,�+�kw�w*/��G�K�` ��"O�Z�zP�$	cq��V���x��d`
�]����]Rfa��LE!Pt=x����Z�/��s��-CI�
n$$�B�� �h,ù>n�u���z�ºJ���	 �v"�!�~6LU��^�͊�%��Z��K_ *T=��b$/x0�0�?�>Kќ����B �M'�T`H����j�SnL��8Hl3_�>�m��7��t
;�a�AdK��}��&�z���C����r��n�Ҝ��{q$��9� �+���\|�
c��ٗ���`�^mG���<ި��"z���Y����N�%�\����>���o�!��?�pZ7�`�ô��wJjn���ܻ�9�UL�X�R��YR�_��:���Pٖ|y ��t}�i������F�xC�����q�'�C�Ca���5|�O��Z ;K<Q9^(1�����T��W��y� +3�e���t���!�1n<�W��Lu��v�!zwl˨���2�����Wq�z��F���3ޙ�� �s�,$f���+ ��(��oj����y�W�	�.��Y���#xw�Q����1�  O�C�;u��tl�(�󭻘�9�co��e�j�T��y��1�	zH5#,��ɡ0�IF|�s�͖�ɗQ^�����r���n��@����o0�j/Rf���;Zb��l�c�|vm�tc`�P\/Ā��]� ��!Ts�\�'A1�� �(�x�S�� n�ѓ�1�?�5�0z/叝�����|���a�X���d����L��f|c�z���8}��������3�ȗ0xL3^�"�m�$�c9F�=�<2
^��5D�eay�I١-�t|M���v���q�Co�z���շ_}�������_��_����o�Ҿ��+G������F���]Z�>5䁕�����__���չ&iԯ}`=O0
��J�7�w>v��|U~�0��P%�g{F�Os�xGK�D������ݮIQst�=�]lί,?�28�e�ш�F�O�v_,<�-N:�̰"5���[��^m����C��aO�۶�a���N���A�5T9rW�-϶���}�6z�®X\ά_�x�Q@uqĽ;����9����E~�3v�J�OB&�� BnYYF�h�R��r�|z	�E@��_g�i��-#?R~p�O��M��o���Z�0��@�ь� F]�	�����6��%$����~0��O��Ԩg��*��{)�1��3UF-u���»:��L��	j�iIl���~�HI�����v��K��� � <����u�L{8��W0��q>�	��a��!�'�D�#҂*��@�,O�v���9��z ?F���e�'V�
��p]֯�?G��,�\���������ǹ�'0��a�q��6�������x%0o)ݺ4��S��t�M2o)���=T�O��G�+��zĸ'˳ꍨ!!e�0�cN���Ӿ���*�J���)#�-bu�ܢ԰���O�\���T8�ed����h'c��i�>��v&��;�T�j�+�k^�����[C?�%F�/eK� C�tU�w�BdBY~����+���4�YC25~^s1�
_�T��i��1ة �efh�?9OO��z�u�%��|�?��nO8��"�ax��.U1��y#YG�ͱ�������R��XF�G/T��H�ϕ��~;�~�$�1�iL�Yܕ�u�X@�g���ZUG��eU'M��? go�o?8��t+v��E�@b���(j��ä�'�.�<Nh����3��gB]���	=�>���}���U�Y�U2������|�)����^4���{��Vo����VVgq�FvD�t��O�:�T`*�&X�G��ʱr��0��LO;U�>I k�Xl��ʕ� ���]pWb���$�ID���Iv�i�h7�C7�U�"�p6�q�w�U�S��Y��F7~�"g���4�rgUݵ1��%j����C��1�y�����9������39��@z�b���|4�Ǘ>��er�G7~��� -���<��q�9|P�kݎ��Oһ�:�{�ʮ���#���B�V��3��/SaǈbdiA�)1z�B�&ܔ��V�6�{��o�d'*���F�&�7b:0�ڦ���akW����F*<�ꋿp�j����6l��ZL����(_�3$�ߩpZ��q,?hߓ��KH^o4\��IY�n�$Ͽ�ɃG�0r ��8+ݎ��uv�?�+��o�h�\�R �_K#�N�-7���"�^��k��L鉹����e��>VР�0g���Y~�)7ZJ`�
��<K�|(����Ȗ��퓻�\�b��d$��ػ��s�m������1h� �T3�F��y��k2�,m䫹ſ8c��r�ȷ���i\��j7 Օ$���n��B�D�[0�s'oIVC�IDH���
���7n�į�ni���շА�K\Bn�E���Z���b"�8����[���[�A�/	�V��;`�U�������ḱt����'Y�b�\w�f(����1m�i&��ލ�(����!�dH몥�[~��	��[C0�*Վ��A��pȚ{7j�<x:��(HHu4'�[fP�~Lz���P0v@;"�2��G�4ǽ��цG-�~�j��F�z���.�ye%�]%�_D-�F�7_�ʸE��d̶j6]�@2*�O{lh��y�\�N�ҝ��R7Z��ep���xu��(�t��e54���@�UK�2A��1����]�	�y���o�^�*��D����9	F�Wj�Ѩ����W���Q�D��T�	��	��8)W� ���;�6�6�
0r��lK��s l�ү���`�x�Mo+��,;��,�ӊ���w��)��]��F|��]�g9�C�+k�J�8�B�jA�Va(c�^`t��>9�5'
(9_}R�|2z�tX�o�Nk�- ����ֽ��{ҧl �`u����ͬۡ.G�^�eȻ�6W����O���7Q .qK��Qi���e���b1�Ϊ�㣖A���������k��I�G��R�I��f�>�l䀉/b[�cG���b�C��O�����}c�]��B�����1y�BW��4��a��~�6';���տ�V%��EMk������pR מ��4�F}�q�v��������/]m|9��55��YD2͎��$IF��������2�Y�VB������n+�%�ro4̑2����)}u%B�"�`���a�P�����mkX�Aއ2�:o}�������@������6e�ŧ�ڻjX��Q��v��ZH�l鮗|'�Y���)79��5|�~RN�%�7����e��Q4���eTȁ�n��F)9��h���!{��^�i>��FE��&w���G���mW�u����R���қ�U�6�v̐�����7Fv cO��M�H&��+c�fA�#���~�J��T���P��ڌ��Q�<�i��1�L
?�u��A�(%��^_����$�q�z���[��&�c�`"�e{�=dp�a
"WZ���z �[H�ߞ=�O��ظN�\v?>��d��<�٩ۏ���#��N�;� �P�:�H!D{�$�Y�HT8JO���	�8�j04�Le^��E�J�<X�c�R�$���޳y5� e�sh�����you;�|��'nr+����;���q�9䭪�<��1��Z�9��a� ��>i��#\�˔��`DR3��&977j@tҫ�k#�*��fk�ֳ�s�_�Go|٫$-h\LwT�	p�yX�{By���v�M��BVw�.�k�� �������_��y=4������u���%������ߊ@�H<^5(�o�2�0��՞�)�ҋa]Y�j�u �&َ����$$�4�Ƨ��[�0	��_&��`hq�xr�M#�z���uO�(��2>=W���U��J����^�<�>B�N`�aV�����W}ѻ]n$4�GG�|.l|��8�s?f���럚eT���SO(US�,Oc����2�FƁ��@��0(��d�ضn���v���u+��B;Y�XQ��	���_��!�!������g� �)����7��<�W���P�h��(�4�<ډ��hz�F7���=�D��eKRӄ�.^&�C��򋻋N��`��矚Qg��*'���׌�1�%��*-�Z�ږ��J��'9���-�1���v���:P֨�:XY�=@CXS�xC4��d�}���1� Ð�����+ulA�Y��J��hEQ2AZYv���l�Id�䞨jF�+ǻ�!#�~)� �ƛ�<M��zK"#�X�2ΠM�t���@�ȣ�Bj*3 ͜�(��p��a�2B_�R\]j�;p&����䟠8r��1MU�?�p��m�dB��)�G0�rn��ܖ��C���C���č�v>9;���v���(�~����٪V9*vE'�D�Q��z ׁ@/4x�B�[���ض��q�@h A����{�Te'Nv�Y5�jΧw�T�A$�q��0��(ޮ�%�3�����+'���b�;n~=�q��$�Ӓ�o�v�[X;rs����E,�Ez,Y��5n����_�|�9J�܄�L��KI�ƍ��HWn�o�U��+��r<���2,!��W:��?�~�d���d�_�jF#��C�� ��B�L�cY�,h�H�������Sɘ�paK9��J�t0��Q,O����]�B����T�|�AېQ�����Sc�)&�:(�{��M��3�!�1*Ȇ�!Z�=�hD��L��gO:���X9[�kS>�Z��XZe>�l�q�l������fR
I_��Q�,N�ș�}y�h4�27>���r�Ʃ|�i�!�Uw�o
jY�@� ��,&��+J>�{)�k�j��xH��Z�ԆN�ذ=�n��!1��˛�Ι؇WJ���ُtw�_qn~�*8X^R�='OXk�0R��>��9���L5��gr�m��d��qzϩS���5Z6�_H���Ĳ�S짙�Tu�z������`BV5�}�tsD�\���Ǩ��o�+�ygl��*�+'#���x�Ǭ��{�|zW��B�ܵ�/3��No\��8�m�\��j5cD1�����f��8y��GhPE��SǗ�Aɘ�~B��͵D��B� ��޴,� 5$&��Q�����֩Ҫ�R����/'@:T�)@N�sc��Z�Sc��-���d-�𙇘0s���c�6ɼ�WS�ސ�÷��Jaȩ�"4�����~�iT������2�G�8W��}�6\�n��}���������r�����t5�Yn���6�F����V�e�VR����`��fRh:�F���1�dxEԓ�f$3yp?kN�n���@SJs�<o���@�����u ٹd��[��WԻ�Q���T�a�P�N1:�u:��t(BT�~gkO�#~����&�2:�XF��Z�Q�����s�o<qaV��#�[�{XtT�<o]��p����⩛x�'���m��<�V�C4��e
)� Ħ��h?=���K��@�$��V��]!�������W���|(@^aR@x>�����%��񫔍�����(����{Y�AW��c��@�	�7 � ���]�a2в����k��-�N�a;����T�5'o�=�9�b�f;�קE%6Fp-��$��]��^O�=kQbֿ�S�������!F�Mû?�Q}���|*���⳨��oW^�(���I�_�w�����V��OƊ����v!�ш���U�9��n+�?���õh�vj�(��=��O_em���Gj�c��/�����܊�(5�zܨ�(�����9/A
�+&�~��w����jK��B-X��Nc��:�W��?�~��"B񄳀db.yi!��coՄ�)@�bp�ċ��ikM��&`9�
�g�͑{J^�'����GG�b+b�w��b���~?�(�E�MY���͓�lm��,������������g�n��NG����^f\���<�#��'��/���J}����礶��+��
�D�,��;qP��rُ�K��'��q�f���	�����ۭ�h�,�Tk;(J�1_��>��U�:n��K���HnH�ZIn�<y�Q Ej�(\F�_�cm��x!����1H�}�n�l�w�7\��n��;��&g������C��8-�[/R�����c\-�p�>��VW�ۡ�[)�hۙ5"�<��JRc}<�R%�B�Pb�~_I��l�Ju 7���LB��4����R�#��T��<f0(I�j�z+��Oj�)�Sm\&������ 9�a;l�H��a�h"�h�l6A�1�$�G¥h�C'�Zw�1J�/Ny�^fZ�es����Wݿ{w�Ġd^��9���ݠ2(á�����;f���Z��C���D����������a%���_M6���%�}��`ղ� *��4�ί7^Q�)j�2� &C.w9���t�F_���J�:��
����k�����bEcs^B�v
5�{<��t�mii��z���?�{�+)nF�7�o�m|T�m���^�𵝴�0�XcZnbe��Q����+D1�AMh	%�
k1���{�˨Tz���rg��<�I<*��)���*g7~�x���<L*���Z�+۔�ڤfU��vSӑ"D1iŊ��;m�3~�W�ӛ!F��~�_��}�\��j=�D����{ݪh,C��蟋]�"xx��}^��#�,�?̵GCNiI��q9QF���uy	]�i��P/55q�O���}�h^U�HXr����c;y�Ս	�4�8�Sw$a>ۂ�ɻ�b@�����?�7'3���AԴ��oǊ����r�Q3>dQ���F����T������lȘ#*z��'� +�J����y���7M�0����-�X9rĠEO�+7����$�����DE'C\ifb4�բG4�w�=}nϕB���>Մ�����^�C��[9�!943
/D�6����r�$����2c"uk�6�<}fv��	
��jX"։�Z{�=lH�9/7 �|H�E�UA��U\��� UjÃW�Ki?n��P��Z�����+f��ԆxN�K����	x/2E,���|��̉�v�о�,v��6+}Fj���4�]t�s�{u�Ǝ8�+�r��`���N4�k���(4}<~=���5k�}f20tjǓ��q�]���c�dyD�N��;r��/M�L0�}?(!`>��1j?�
̉!8/�G�p:˝o��v��U�A?�3"��x�!�(�)�ۊֶ"� ��[�0eg�_���-���R9,�"p�X� ®��͍���y����oW��؏Yڲ��?��+�5���@���;��l{�R�y���8���,@��0��@B�;-��_��b(��J�'������;�����J/�ڔ�#ϻ]�}��b�͛6������~� v���Tҗv�':/ X��֭l����;��n�1P����>PX��UMj�%lK%�%��.@�H����"ۜoDxF=��a/�
����tNT9�ݺI�E�?�t[��aɬ���R.Ʊ8��s}}���k.�>`���>wdW/��M��H�̹��V㎅�4��
	�,��Qv>j�M/������e�����ix%��uy���ǎW锂
ĸN�CD��R����{�O�P��H7=/7���O>���&�֨�+*
��{�4��iQo��b9@�4'��Z|�4{�H��iv�������A�n����>i�v�Q�y��({0��t�3B`����A��x�	�G�8��N,�$ �@Zb�!F<X^�O%���ԍ̄\�>X�����W��ʬݼ���L�u�g~k�|��3�
�S1s@h�\2?����)���cU:�^yy��lA���dV�kj��<zs����x�I���,#�@'�(�f�hF����L���p�79E��k���@���?��lF��d�z�a7^�5�F�fB�n�I+R��ҭWn����z���hi�F ����
�?�D��~.�g=����}n�ԅ�fۮ�
��)�EkN�Wo:��آ��o��ȑ���Xh?�U N�XӬ,O6c�=>�&b��,=W���{�T��#E��:��5���˰�&*�jxP��:0�g��%��2�ޗ�S3"̰�\�|���#I@m�)�;F(��83#�b��Z�-�G7aLF�XV:���)��v�ތL[�<D�c7���^����<{-�-�{����S���Ճ�@�I��sxfƘP�
�2KHmf�&u2;��)C_��-���#ݶu�o��?��Kvy�=(>Ɠ�-u 傕�]Ξr�3o4��]�hL?�n�ퟕaP?�{5�Y}�9�߲v#��/����g�٫�qO��E�x%�_Ց�����B�]Uv�����t������;3|*ŏ�樑�G��9d�O/�_��ͭ_��=�LBdd�Z�k'��9�լ�\�9�ň��w@���r�c
̙����+U����IFw��K�v�v^�����
v��5t���/~p��_j\I�75���&����`�D����2:����\8� �u8M5�nB��Ix8|�Y���P�I���ثw�d�E��E:l���Ϸ^�P^�h��φl>A�[ ˛O
Pc���0�������Wڑd[���^�ɨY�K1\�����0�Hm_;*�=��Ԉ���U�v��OO��
G��ː^9�̐\w�ۮv��y�NUp&�A����Qu���Ʒ��������UB�lK�u���#=`�#4���95��e8�|3~'v'5�x_�|)� qUv}��^��qQ/��#�je��g��ވ�@����bJ�5b_�-�FS'���3$v"Gr�nq��ה�R�����xL�*!8'��v���^��A(��'M�"y�\C�k��"��RVc�,5�x��4X�[W�^�q~j�� :�=(�nG���>ܴuu�z���l!y�lH���Gi��_ /R��*���'���uU�%�4P1��T%Tu �m���Y��73&i������<��)R�2Q>[ֲ?�W�坨��4�G�S�芖8�[ci�7�=}g�</O�Y�;7�u��U��q4�鲼���33�G������vo�8��Q}��$5|0�}�:!�G���>�lg�^<64c���A�m�)Y�	od�x�U(Tй���ѥ��䫒I�Ɗ����/w*�d(�U�~��K��>�K?)-8�Xj��P����9^���YyDsc,7GwEy�+Ɲ��9��\��� O!x�0�^�����D��@F����l�o���\�̃���6O0�F4i_:^%W��n�X�#��>9�~*SG"�XƸQ��ah�Ȅ�7G=�'7�L��9)��Ș�ЦM+G�E=��ba��Y&�mΧ��I�Lo��Z������iֻ��l�!�i:��{��$;�A��G��a�H�lMZ]	~Ӎ���bk.,%ͤ��/r>^��qܕ1�=�GW��|�B�u�n��#���zEmR%Z��B\(���rN�R�����ϗ5ͩ��_=��U�� �8�'m��h=������̫#�z���Db�D��8T rb���j�K����N?![?���b��Rh4�O?o�Tdq?�h��P(�V�ԍ����ʡ}�N�w�h0b!�>�DMG�����A2�Llc�iE�[tz׈��;��\����u���"�i<*��.j�����Բx�wV~��	���5K���x�BظG�yy�2ݨE:�'jST�H�ۃȖQ�鰶b՟o�P�,f5�:���>�n�Y���~+r]=S:����!���a���������T��F��3ٍ��g,��o*::�o�3b8�+�\�͈2���'!)嘒,op�b�	�Ǖ�O6 ������.g�Pm�*h��?~�4�y�hc׬2(T�|ҀUΗEkY-� 9���?�Ċ�[�(�1^m\ Hᮭ�cVS�oZ�~�`398�A��{�v��z�#']�8���'(a��Z�f�S�P�Tw��D/���t[��kǽ�ń4(�+4rH������j$�+UU�Zb���'m����m��)E�3_!�l&�s��=A������;��'�; $}�Z�����9C ����+�@qI�=�+u[�M�.���x�2�T�L�7�D�o������¨�^?mVW٫���(���I�$d��E�w#�k0�����Z����V�T��1?������Bڰۑ�]�!���;Z��n���������oj��+U��۠_���WPai=V=�kXDz�|��!��H��3!;�"�<�*����2H�J� ��o��w��P�~�oj�R"�֭� sj�ߧ4���?B$�?��L� Q�ո�Ο
HR�~�iu�˯^b8��S���$�+k�
43�.�6am|1�6��Dy�[�Am{�*�WF`�MT\ft1��J�!�{���	�q�i���O!K]P����4�<1Z� 	(%= ��"27�%�M�"%&�S��p������s�ܑ��1B1O-��KKTk9�~���Klc���LU!̧/Y�o�퍍�P�+��Q%#ϛ�NVU�\�pG��$4���v����r.m�f�Ԕ��[�KoO�7�U=�h��8��*J�����*�F#ga;>��x��^�Ч!1W�{'8xZ��J�g��l�tzg2�14R��(!6e*�٨w�����h����Uey�����j��3.�2GПԚ�3։/XVK'ͯZ��sٛ�l�f�k��,sE3��F����٠�|{��|�[�c��
�d��y<�pr���d.����x�|X��;��GΤ6F�v�p�,X<��l�A�5��/�/0���Yo�JWV
z��8n^�}�ǜ�ңۅ�!�z>��͸sT�y^]��j�"[2I3�䤦.Cd^��{*�lvȇ�A>�0'�=�L�>G$,�'VD����pԷ~�iT��-De�^uZ��}C�k�\��QG"͘��q�{S��5��O�h�D.s�*�n�,qI�u�&�9@�PIq���S'�l�^��`=͂�B(�Ca҂���=(?raOB�}�`��WH���Ygd�%K^��X=b�]�}�^��гzT�R��D7���M��+�O^��Z�-��h�D�uܝ�P��V��iY�� �}�e|l�U�5,����B�����$+�z��aί�I���k��{f�Y#�r�a����]��d2�$K�QR}�C���Ɯ$�ht'�g��8L�����b�J{�U����KDft=71쨵e�F�"���ԥ�{�)W-ԽS����-�P�ɼ7�Z0��XX,l�癬��}e�7��5_%��28[M�^1�H��@UU��i���2 ����21>��Ȉc����fh��)	{q̯��@�~���E�rZQ��^�Ȧ�}Y��*�v�4�����%���R�#-�I/�Q:��;�lS�n;}����%�k��W.{�c�7}?n�Z�;��'�q�N��#?�����5R��{~�~m�� k�I��[py�_�O��uK}���Qj�.t�ￗ�pZ�S���-���B��/��B��/��B��������oRRߒ� ���B������S�J��
1�.����ߌ��v���p�c�OJi���no����5Z���.5Գ(_<�>�V�xO3rc��`žK���酱��^���>��b��ӧR��㗖�II]�i1�zG�(R)��MMbo������B��/��B��nΉ
&�#K��=�I!ӛM���������Fj~~��y�*�P��V�pc��=�_d��vg��#�S���ۤj?������x�tU�[vm`�z�\�h�)^�9p������K�Z��2!y�I2�g�e%s��yL2�%ɜ/>����_|!���_|!����fCOwJ}��ڴ�e���k|+�f�z������x!c�t#������w֝mj|\�,�,��������K��PK   �A�X�l��A Ԥ /   images/670050b8-4f2c-4603-900e-28b8075f4ca8.png�y8�k�7~��]	��%KE�N������C�Ⱦ�R�ꤐ=YZ���Rq�P��/��/�ݘ�����8�������/�u�j���z��g��Z��2�1 Xگ�� X���+�=j���U���� ��G��ϓ:��uW���cs��9�����I�OkK{�s��m��"��� � �W9�9�"ul�Y.�Ov�V�Z�d$�ί*H:�y���Ե;�_o�њ���>ض���)s{��c?�������?�#?^ia� ��Y[[��/ﮫ�ŵFFFÞD�L��gF�O�w���}I{�^�w��+���v�^3�Rj��o �зov{�������ϴG�&���*��z���E�]?N�z�Ff[2�3�͂\�$Y�\�p��v��NL�
�U�aT��?i0�&��}`���յ)��Dt�� GGG�Ș_�ҭ���y�8�X_U�hʫl?�7Bt�$�Mр�o���)+�2����G?4����%G�s�
'򟌌��?98Z�	zÆWt�	�����kk�s�r������J�ok����v�v�G6{9�ى�Ze�Vf�ޭ'��F�L�����hϴn�O����2S�'i&ȣG���"�(�i�4�"��9;�����R��Ӏ-��~�],BEF�̔�X�X��H`����Ư���{j�-ó��5
OW|]���YH����dm�j�~��uW�Y�Ke���x@�
.̒��Ʈ�����&f�&��Y����{��'F
�R����Gq�۷o�V����IƓ�Ñ��2~��b�y�D�F
�Z񚠃�UVK�&(v�_���~�M�7��~�M�7��~�M�7����0�y1��?�v�$�g�+��[�r�������D�=��DlM�ph֒H���\�����+xJ���?j���ܼὓ��?8�*D�I��x}�eT�ī�~y'Wk����H��}���G[Z�?1�7��o �fZ�/yQ��/�~���_����������T���0!ʩm�}�gf�a��R�k��ƍE���]R�)���Q �i�K� ��]o�+�+x
a&���Z��^�4X]���1d�*-Ԍ�ʳK�h7���Qu
�mKdLIG�("|�n�sj�����R��~�9[)ܞ辟��?_�-tx��e?�t?a�]�ȉD�a)� x�`�K��S��'�������1Kl�|�����aHnj� (�I����dN�g�}�R�U�e��{���?B>��м���zJ���2�g��Ϥ��!�B���sfU���Ś�c�x�����C��]kH��!���G;F\�@�Ȇa���\���{o��++{�,�C�R;I�[Ӊ��2�y��b�N��L�/�J���άV�^[Jzs����f�+y��>Ȓ�m������/m/��WFF����1��'pU)L��f�U�SJ�bH�e �NM�w��U<":��D����"!)K�.e��S0�d�-�EBD$!䋩�ܙ��H�1�e�3�� Ğ�����T-�݁��ޅ����֞�Jߎ �����!&Bk��R����qШ�9�*vU54���k�F�+!�4�A�Wv%*}N2$h�^WY ��E��e��Iņ��i����îb:]hNJ)�-��G�g[H��g @�'ݽ{�8裇&?S���V��̸1�@J�e�R�4v!XBt��1���4/ba�c��P�_q�8��J�ӡ֢t�M��`�����J{'�荘 ?�; &�OW[K /Q[	�pw��Z��Qi]���>k|�->��q��Er�| Џ�I@,��5Dn�IêI������"����e*򊮘(��>\�L+of$�M�2U�儐6g�@��t� �o{�*� ���X�W)�.�'l�GA鐪-��1bO;��`�I>��&?��,F�w������ߐȤ.�F��!*V��t0�L��|)�q�`� k>�'xM;�h�� F���q�Z�n_�����)H�+�v!ZOr8�7���	e^�4^��:k=]B�77�a2�j�_e ��/���+��[�x���51��-�.=�{6~I�(r)�,
�+vv��(E|�,�Ξo�^7;��QqQ�P���2?�]/9ޥ�[]ʗO�˼s:Eq�!�t3j����I���G�Κ�M�P ����O�cn~<65�*0R0e�?��6F�a'�[/�g؁���<�4��3��1
.S�N%�B^�*%"Ih�$��%ݶ;G��&��=��T��V��q�Kz߸Rav�٤���F3�%O�֒�/���K+��I�+���[s'T5��D�0s��QKc &�ۃoi�z4�Z�5���&�a��He���MQ�QF<a\{>��n��F�]���os�їbƿɗ'���?�e���t"�"�aAP$�H���6�ᢍ_�0#�2a�k�'��V0fm���	l���	�"c<��,�|���c�5%짞]	@���;�����k
��4,���1���z}���Lv6p����J��+M�5�C�E����NYJ���1et�r���7� Ds�خfO���Y��"���*hsq���/r��ɿ
&��b���o�H�W��5�����l��8 ��A2o�+��u�T���e�;p���b���|�zP͆h�Q1�d���w�y�I�?Vp_�i��^uV��EЁ&F[�A�fs���ҷՄ��oM����B7G� 4r��eZ�^%���?~��x���� Æ���a���φ��g�[C˜�5<�֭�F8�*w�/��nt����n��-n$�1�{Z{*�[�My��u|�K��*[��.��"�N�	�GBI��z�Ma0��t���).�u+�="���B1�d�ǬO��1��u����҉8P�(K���DV�Q����K�3�'vS,fpW`T��j�v���pފ�`CǙ��W�p�^���X�U_<��ƙZ�K4�*��l�CTe��\�
��WAJ�#�A������)-�6�"L{���}���F���M�0��`�d�j���pb	_�v�jI$�%�f��O�'��gmN��~鄦���~���fq�\�iħ�]؋.�o٠�aPT��\�� �d�������W���WV�X�mԽRz.S/'��m�(0~o��;ݟ1糖���9��SbdBH�iz��	��4�a���/q��5�c�@ ̾��CFkb��d�;��ix�aY�#�Y[�ji�ih�yC&���/���HH�q��'�a)�RV{��#�r�U�O����ceo��$�q딃$�6����l�8op��9�>�T�b�vI�������M�N���U�J:v-2�~%0����o�} P�Zt|��.�_:`���+��?����?�%� Vi���\�cz�k��\�K9=��9�a<�O���X�D�!3�ь����P6E��Z���xLo��&�a�C8ı�}{�J�@�`�4�)7��J��7k�e��%�ך	#-���`|0��6a7�׿F_�۪L���\�NN-\��#)��;6���H	���m����.�*��U�D�R�2��)�B$q%:�a��>�ХN������!�����d�{?R],���~1��	���Zv�k����Y1P�C�9�Ֆ2��^��`>��g1�<�Ki)�VC��c��px�p��5q�F��̽maJf�����x��\Z͖W#�����O�১;����A~�
��Q���l.�Z��̮���(�t��%�u�y%��2x���E��+My�'�����
����o�V`F4�ݹ�?� �(���XVd�]/rS�����ۧ�0x�#A�{2��J:r��~\y��_��.��X�ש/��I'�d��1��j�Hx�UVnZxV�?�Ue�b4�l@!O��z�?���C���3�B�g��p�'�T�Ӎ�y��o<�Ѹ�1��`9�q��|\��znQ�񯑦�Ƣ	v
��]��D=*�2a�C�x�[ͿGK��^qD����.�lױ�ֻ�����)J��|�QFy�_Qv��,��(��ϥ�H} �`H�(��th\���1B#�wV��0
<��:�nE�e��պE��0��ԭ[u����T⴬~�z;��9��c��K��$���u6#���?^��L��XO���O�JY39$z�r@�e��&�W7�+��]uV�UJ^���R����T¤�Wz�+����ldU����]�ݪtə�XѬT1���93G|�].0ʃ��jg���ү){K�=$�*��r?�G�k�ǒ����>�4��YÊ��4�JX� �$���rn�8��4K0���e'�͇d4�Ϡ��
b͐Y6����u�����/��0�i��?5�3� �oL��Z#�@~��q��l�T��Ɗ��Y��V�ϵ/��.�-ҿ���K2�Cɀ%����b�
�7���;���Dҁ^�P(��a�����sf�1��_M�,xH�
z��]�xl�� GJ)W�n���pkީ��EGC��?>>O��ű�J;�VW��w6u?��T�{��'��l9��_�{�Mn�6>�st!��,rȽ}��%����vb�G&��9���ʘ��7o`7�W�3[鰼QJ��Ӟ�!��q��GmLj�[r�]�8��H��H��� k&<��[)Ɛ^��M�?b�Co�;��e��=v�HWF��ŝ�V:Ac.z�x���J�]��|�1�;���K,%�,����6g�>$����x��y[{6�����t^D��ύ��6��
����A����U�'�6� ���.����n�wGb��ۉ5�xV:[�P�±�)u\�ݮ*�5{�[�%[	sdφ-여4D	r���g߅��*�OWKe�DCW�W5�`�)�ƴ��C��s�ó;�2�����Jp�㽻;���H���#N�t�: �����VZId�+�)U�H���k39�����"*##�X�Nh��`+6�i�/:��<8�y�-�$�CqyL��l�rl����o������X��^'����t7���e�����3��[	�F��r�p�U��3!�m�5���V ӱ��_�c�W쎬�*��7�c6��}yt2NHr�o܈�W 8��T�����N�\,��e�6��/�_����穥� ���E���6�| yY[�}��]%�y)�u�#/��`�)�r��U�W\�>lA��y}0���S���D�A�Lv �G�F	���u�J7�6�.�xm��l�\9��7D������O#�؍�����E�N#�i[i%��t��".Α��I�92	+�c=�!�C�0�Z��K�O���$m�����l|�r�G&#��ΣBt��	,Ƽ��1�./'f=g�^�i
�`�	@�a��hBQ��'����Ei�v��8fvM�<�"�s���3�Q̺�'~���O°Z�<��ԋS�
͙f�S[n]T]UTe���1SUU���h�W�3������o��gRpo�j�����<�{�[vb�9�%�^s�,����Lc'S�%�"cBA�v�%�49c�Cy�Μ�샏g�<45���1���
{�k��L淶G!Y)ݭ�8�m�3�nS�QS��3O+�m��*�0��9�{c�&��KJ��.2�H�܅�f�9-;sD���SB���tP�����{I���F3���t�P�),�����q��rT�Jw����~�$I���ْ8�?�b�d"��$)N<�3d�`��`�l�ia�w�ǅ��,�>K]�'�<
YX�0�;�j:4�A5���X���]�)�\�DeN��:���H�t�U��҂��<=���x�tz�}����hX G�ݠX�k���D�u�}o!w���Y�^����ʼ����d�+e:c�U蘣��F�2x�@f�(��m�^��EZ}ѥ�y�`atOX���Ң$����X8!�t�2�&l+D����28P|�f���s]ܹ�E�o[h�mY�@U*�߻�Zm.��5v���r�r`�	���9����9��2Zݷ_^ѣ{��lC��;c��c-��M��̗�.^4��e��ga�[��[��I9U<�eCd ȧ����G�;P3�?�f�}D��bb}'�h6���V�c��i�#�
e����3 6d�N���M?w��r����~����~�\���~��̒~��I����[����J�cѪ,�SѢN ��M��W'Y������"���@O�04^̼)#F|��	��\�'���*�d���f�p�b��da�bv��;j���-թV�� }X�N.P'�[?.�^'��#u*S�2���up�����q�Ξ'�����p���� BiT��R��"@*�����П����Ⱥ�YÓ|K��cA���,4 H�d���R���ێ�"��uq2C7>�����i�ԁ��p�)�t������+T�SKŗ���0�E���*?��,���[�z���_�m��!RB�,}�|Ϻ��<��F�}��l�2S2߬���GY��0��n�I��ʼ�>`d��g&_����n���g�brX������8t�`�p�R���V�o�L0Cë^�����-H�l�_�'�_ލ�,���xB;<r�\݂23�CW�~�z�s�K��潄�y�jŉd24&���Q�nȐJ�K���u{a�����g��xhc�����p�Ɔ��[<qn�C��T�����@M�r?n�:���&�{,�5oV1������[O�S2�	�E!�;fDX.�9���v�kh�ِ�ꛭ���g6t.үo5�U�ɻ���N�t��e�A
Y� ����:�*Է��qt�F`���{r0����HI����̄�V�/E�{;ȋBc"�I i�BԍrA}�[�������#����{[o�ԉMx�ÿ
��>�_V��E���V��}T���V
���eӰ�h�!�r8e�F�A+($m�� hN��B��U�W��(>B��x��E!�^��=��g��.-�F	h�r	���FY{A�.ǻp[���Ӽ�D�r}���������݃MM��ͷɛ��� -��'�,���z�u�Q�HMYZha�!kD>!�lI�#�U� H�5�i�8������	���o��Յ)�,hD6��Ɣ���q�� 7�K��k"w�����Nns�\U=��9�m�%�~Pn��7��[.���{#2���fr�G!��[��$ļ�v��1#i�{���/��< �Z 3y3epuj�uFn$W4��?�e֓8�:����&)�T�?uɗ*Ll*�����XG���?��T�ݼ;���b9?���塈���n/��)P�,���a��$��K`F�
�pJJ��)`w��PsL�,FQ�s��Q����#��co���J�o��px���vRe53�IԈ�W%T%����9��h@Gr��qDc��b-������aff� !����?$j8�%���xA����A�\�l���7V��ei�)͢��m�Π=��s��_�e�,�7��oQE��fV�q& al �"NND̦�=��6�<�3kzݓ�&dץ�|e�A���/��L}�t�
s��D��'�>��=1%��s���;��Y�J4�yD���6g�DF�}���J^<0��Y��t݈Ԉ��������O8p��CWi`�G©@y�v�%,���$�u�X�?cH����p
��� p��)�Y��\0�ߖ!�����3fo9fс�rH�}�" �>����Q�'�$�π	�5w�g[㰠x7���u��R"��%�/�m�q�gVK��[�B���(�)?/ ]��©�8�j/��$��2 �i�č�VF�����e����(�2�z���$���/���5�sٿ�ҥ� IC|(�^�?�l�������Ֆ �|#Z�����QGD�]Y�ls�Y�bp?NNY�?��� lފ���D!h��q#���^ |[�D"Dp�y��̼T�I=#l���M�X�6a�ƍ	��o�h��6CJw"��}�!���e��j���]��|�*�F�Kt{*tI�$O�oX}���3w��722��y�����o�{at���ϛ9Î�|�8�Cx��F�O�.l	�1�p��M�E��,��ӻJ�c�uu&���������fg�x��%� :��$o�x�����9Xa& ������;�yh��s��/:1��<�E�%{���_��eMn�w�'1 +-H�Y�KO�*c�xh�����M]��y�}N>V��8����\Hs� fq��>���>�,eee��[1�]�$��I3����pW���Sp^s��ٹ��s�Fj�,G�.h�L'T*L6UFi�r$�8�T�����<vB��bf*B۝�CKf�M�h��s��e'3e	(V�e&��J�|���2�/GI�/Gt!��Km��m�2��х8��z���sҊ$�n�0:\�zc�|���р+���g��*���:�f��43�\�Hܸ�`0�Scbη�|ĘE��0全�h����Ħ
g$Ұ#�R�[|F�9J�x��x��Gq�U���͆�YI�M�gj,]N������H�wT�?��P����Z�ј]�]1a|&>>�ݍ8�S���4z�۫���\(X��5Ki��z_�h��֋�s�����R����>�nz"�qFM�4����K���=�E=�J�o�@��?��{�Y�������l�t��fMnI�xû4�'!p^v�eϫX]�p��\��ff�h���w�oy����;ٔ�N?��y�k_񙹗�yH����q{�v�� �����\���B4�.so��|�#wދ�=�����˵��Zt�r S����3���uʥG\.м����p���hMr��I��ļ��αܻ���;\�A����.�$�q�z����b.�$��րd�*�Z�?i��$<���V1TWwv���M�m��/���O0���K੖�n2��|�U����_���k�XB�C���[���=tf3��C�l��t���:D� 8v@���z�SQ�3Y!�Px�ο
�w`�~`���N���J9�h���U��t��n]�p��m���sݞd�pd,�#���ݕ,U.�ߟ�>���$@sh<���T=3.{�o��@�I޴�g�h��SLc�ǣI�(z� ��VB��Á+���/k{.��І�j���.?uNa�=�3N�W��t���γţ�f]��f��hb5 W���ڜ�GH���xպ/��QM����)Tg���D!��&��\K*
�Qz���
m�yg��4�U��'�$\�6�iݓ����)wgC�K��;��{[�/�:m>Ro��GE�^����Ar�_�����Eu�V:����o؞ڸp 0K_�F��i��h���=(�S�,�[�u���E�W�X?��I�� T��ٔ��%���H�Z��,s>�����J��\�]��; �>�<
9f!;�8nv������N�Wu�!vr�}u�{�^��V���DC��^�ɯ?h*����B"��{Ty�h6[��^����Pa��1�<ym,?���ڌb���K���\JV8 OI�gVx�!v��b�H"����=�<u��j�"������]���5V�oh��My��ho%�B&H�~��:�$ʻ��`���q��~R���[C����n��ڂ�jP����	^��V�D�(b�M�}+�������2�F7������8Wfhr;�"'����۞�WR���Xh�QZ0A�r[{��t���1G?�!uv�}Y��: _i!��T�EB����t��ޘ�Eά��q��;�I(��[�t]��-T�L����S
^��[8�޼v�B/�,��7���?Y���B���	97�B8`��$A=�\)1��@�����+MJu[J]@�*��d}:P�P��^���V=���B&��54�n��M�[W�O[�'�V�g�Q�U���N��A�5^׷j���GԼ ��2�v�2�+��x��WvI�Z��2]�yJ-b��H��S���ș[�����ul���`^��е7����_��Ey�TC��&6���1s���EL�wo�D�tG�"�Y�r��k(�@�dd�p��1�o��=c<� D��]:E`f6J�k�)�QRqZ��Q)m��Ff�G\\rS���>G�!#��_�[�R�-��.m��/�:e�J�qs�`$QN4�_]�u����=ֺ>{UJg����bC���́��!�a^s߾�m��U��I��r+�E�s���O��ObHX�L��wr�H���!��R�^���`=0Ie˭{�KA���s��rb��W�)�6��<��`���8S�X�����ɔx�gY���"��a�')�X���J+F�V\B4�5�A�	Y��"Sχ��#豗`;�:QK
@��z_�kl0E`�MX����&?&��4r7qD�>�d�������> I9$�?�I�	����A��0+�K�����҃�qRL��`ՄoɆ)�� Ƀ�Nru��ky���8m��	��A)�ܑ��˥��!uR9�&  D��OM�q�tq��a:�8�a�B>�Tu�c,���`��ST:�T����ME%ϭ��銟!��ϋ�^�B��	/��y�ۮ&�-�a~ɷ4v�K}�Ur����:V��C�җ<�`� �I�j���P�;����Vw�߸�"+�����(�#�CH��	WV�}e����˭���X?���~��~��_`�P�3A�|���q�����r
P �����2�W�a�q�҅��en.�[wi����v�:Q�G�{�N��w:�H�%zF�T)�(9w����|dfff|Lt��T�T�n~v"#�`��"N_ܖj��M@4A�U�p�����d��Z�%��A<��)$($d\t��T�h��fG��s�����R��쀰��N L�<�>�J���w��X������C�}�3�9$�:��ۥL��:�-A��Q���!>�-Wi�j�e7�Ub��o��7�������}͢uan}*X�[R��{H�7ܥ�ԇ���\]gu�}��Vb��
6�����oz�'N�U������sH����7v���R	���8���͢	1.C�XO�'+�Vt�c�,{��q%~��{�.C}�j��*yB
E�
��0
��{�z��1qW�x�۷O;�{���-�d�.���Pe�����f�|nv�(�G�y��#� ��x�)� �k��	;� ���[SSS$3!¢!�8L	��� @��0�`LK�����yj�>'v`��9T��Ӻ�H�@���uv�܅��4>(�#��Vp��Z�*��\� 'K2��� ����W��I^�>�
4(���� �Ox���ЃD��>y�
���=��4�B^��C��(h-�Vv.�^������(wikd�2
����d�8Q�L����J��A��&<�������,~	?��Y����t؊&H�A�&r&o�v�4 ����H �?av囪�9��g4������H���H�.��a{Z�1Q��!4�ˏӴ���l��R���D���4��*a�+�>��]M3��6꤮��	s/c�lmR�m��n9��>�h^kck��l
L�/�@��́��f�$L8��.�r�~�X6��c,��:��<h'N�x��/0v��ܢ��L�<U��IU���#;h�M��ɉ98�͜�ҡ���U�QQ��I��ww�z=�SHq�">��}&pO��h��U����a̍�K�-/F����`B|G�QASk�� �*���s��A����Ș��M �bB!���h�����:�������\l��'��	���0ӑ��z1=�\|�x�4f?�6�	��HU�	5Cc6�5eZ��g�&f����Η��/dZ�[��t����"T3�t�'|���R�G��q=�{��ɼp�| 9j��(y']:��؉M��oC_�<,�D��.��<��*�K��6󫌳��:����p��1WC��k �ҭ�XPa�3�0�ј�'�C�F��A8ȚIx4�.4��5[���Bۿ3�r��qG��s�1{H�C4��?�L��oӷ�:�4h���z������������;w^Г{A�R��#�Z	��s��kj��+���l�q1��t 7q8vE,��V�(�Rl���b��Q2��K�ǿ�架]��0�4����l�r�:��j�^Pf��c�=Q ��ΜK�p�_�5���A�2�Rl������D"����GϮ�&u�&��Q]4�BB���Ք7��ڏs`��!V�a�&Ѝ��{��;~�=|5�|��d5��<�����L�x�W�5^���>�L�)e�;G�	�h//�wy�Ш�
��O쉾��ʙ���^���3�o�aT��z�rM�d��s�,��hdE�����?�է�Z�#�n"WJI_o�1*Z�3�f�q|m��-O���^z�G��oJ^��D��꼺�wT7Rt
3_[6�GC!�N��VuH's�׈Dq:2�u�H�}P�x��ڽ�g���1�A�4D���t�o��qΈ�p0��F�#������l*��3g8h�kC�2yK[X��Dm�T�{�x�V�O��{�Ֆ���GaM|$Q�M�A�rL:��
�%! ���{9ƪR�[���,�|ӟ��XN�&�><#%p�����,�	��5y�oW���nt�/Tێ���]1��z�Ldyv�1��lja�D��q�
��b��Z��|N�0��,�qe��BL�jЀs�ۺ�-�"��R��A�W![� �q�Ar}����x��:=ݱ�W��h���O�D/��ѡm�
��R6��vX��mˠ	�FB㞀�۲�dh^L�����-�����j�t$"f,�%��.Zr��ZH��ֿ�U�+���,@��^��4�H>�˭G����"=pY�m��b�,�(\��,2��f�u��)�S����ƺMٻp�a\-�*ք�<�ů�����I%{����b�-4�n��2�{ ����P9��y�������M\^*d����ɉ��!$�������p�����rك�R��Ә܅V|M5̎�#Ǳi�R��!�����g��~8�W<~.�x<	�>�;�/��k=h��ভ��!1o���=G�C�	���2��ˍ��/���c+���9j#�����:N�i%�+d{O��r��Vy
�=�VGV*ɣ�Q��SZIFD�1�2y��M���:�� �ᾦG>�|� �'�M�']���U
������K�:1�FY&'z-��*3������0�9���-��� J�;ixQ���oM%%nF�� �}E�/�L?
�,Mo"q�u�r�u�X�(��qS	�dH�"��n���q�������ST;���AU�0q���:V��P�"кb�C�}p5���h���X]D"�!T��7��5�i����{C!T�zQ�*��<B�|�$\ѝԞe]�MY�ӘG P/_�:
�#Z�Z��W�a\)�@����5�v¸:\���q}'����&9�ڐ�ut���6�FH���m�ز=������0�4X��*he�!:w�*u��ixэR!����������F ̿rj�)N�8�㍑ST�,k��a��>r����5����w���J
��Fo집�ǂ�Fߤ��ce'�[ƽuSfxL��'�C>�����mA��z7O0���K� Ǯ[N[C�Ou�GI��O��� ��gp�(1�tuu���?�YQ|:a�x	��|��lN�gcva�H�}=e����@YYY�sWi�R������+��������M�#���v�@�`D�Z(���".��eDR��RM"qFљ���.��̪��*���:��L�n3����#����]{l�[��W�x��+����;��A<�
�d+߫Z4�j�ꩴk��G���4L���qw�L}g]���c��
E9s�U��C!���'�,�����/��+�󘚚8zn�����H~���2�BfM\OW��/fP�~�f̌s�,�Hb��.?�)�`���`x,g3����j,��H��٢��E��ˤ�ǐ7N���;�����u�+=О��  ΃%P/�WN V"k+US��B_�S֗Q�{�K*�9Bc�����׎�r'?�0W �ǵ5$
�gr�_��v0�z�ZBc%�J�r��g�j�Q_9���#�����`+�ty$ڕ��vN&��/v �����S�6d�� 80��"�Oz��P�X���;��.|�����x��b}��n%�"���k"U*�Iy1&��2�0[#g��f+��������b�4��L+�F�ݭ0Q���.��q>`M����iF�J��{��I!�R��4��ݳ���31��J4`쉐W�k�c��pC7 )�E[g���J�5s��#���"�㔶�B�8��t4��\�=B�������]U��#�>�9��d�*���K��^��|p�p�n o��ID'�W��w�}Fr�#2���*݄,��Y����*M%R����\�Mh�6K5�ט��&|��Q��s�C��I�5�ū���MrM�L�Y!�t�M>�pc�g��	Z .��s=���^���v�O��ק�q�N�p��V)��O�z�����`���zPzjb� �NƸ g��om'�Ok��������h���}<&�T�=����"7�<k%�ۂ��a������R`�1S��!�k:������}�Ki��G��y��r�ouk*������g��,\2�p쪌�ښ3Ԟ<*Ο��V|}c��4@)g�j�p ,!X�O�xjLo�������g�I%����fL�0u��\�
M�u�L�ޑ��?;�5������VM1�D�G!YF�`9d��q�$�ɫ"F��k�cM`{x�X.��J����}�\a�J�z_����h�*�b"��e��T��u\�c��S�q(�������v:[c(Q�m���m�+�nk��^('���[��((�-v���e���_эr/�7��A~��Ԫ@����#C�AR�\[:<�rd���إ���E#�>2�P�ïm������pgfؼOe8d[�#�.�zB��B����sXh�2GϹ/4�'��]��l`�!����)�|1�y�܎��"��4o�@*��3��p��Ek��Gp�N�/7��6���C���[n��?S��� ���ɻ����9w�����@tƹf�n>v/eo��a"�8J}L~��d5./���X��TOؕ5�:;���������/��M�G��p!˴��q1���҆��a�k����9�����OVo,-��>ϗk��֓W�������g�h�i��E�8-W�S�S	���TE���<;*�A h���?�H�V9���H���M:B#:UJ	!�	Ӈ�pt�$�b������/���6+��]8�ñ܊��>ytI�A�S����hv���@�U��r7P��5�
�УZ�c�BѼ���r��������,���7�f�*r��-�������`�=�T��{������'��.�YP�i"CY�Y����+G*�3�}'@Z4�dR��$rL4�^|�3)��u,+�R�փ@p���,�3�9�a%:v��bO߶�vN����i�c���ȼ��[;����+�"���y2+�71��d=Bm�?\��v��v�~��r�3��̈́��Y-����:H�l/��[{�:˪�Cg��@Rt�~�Mp�惙�\_'�f!�f$��C�IA��i���E�i~�+Hfd�7ft�B��:��=���ކq��P��J%�D��!祎�\�~��F�\���@���x.��ذ�]���o�7/,�3�xu�bFձ?����N����*�(�հ��0��:T˟A5�S1�OMW�wPծ��=:s!��v�P;kʁ������!Q�8Vo�(�x�d�C�X���\XX칋�	ӟ���f���){SeiJ�Y���oȞǠt�� -��Lj��O7JS8M+0�p�~��]��t>e�Q6�0Ԙ[��|�I	� �:��C/��.�Q*u��ϵ|w��#�n�������+���u���� �J��~=�\Y���M睨���lǼ�v�6���g�ܥR-���vR�k�PI��]L�|K�=�`�e|�$�'�������H�����Ut��v@���?K���.�K���J�~-jP;�ݪP���<����,Y;u�ݧ�T��	!��	�%u|	jױ�]6Y�`:��P;:���AI%��%
�����ub-)X��{4�Ïeu����^+x*����2B@Cn���İ��n�D��D�*�� �Z���B��7�[=��������uS�Γ�$�6�#���T|��O���A��V�?��֩�.�#�6�������o3-�Fmf��άt�"e�z��+|q
J}����,����I%���?(cPu$y���z���>Ք9N�vW^i�b���B���jx�3�����ڱ���f�M��iIA�Z����o����-�Zd��ǭ��s�y��Ǝ��awf�m�?��m߇{)#�%��G~�K�1�&�/��}����}���$�Zr���μ���uB�����KJ���������%�jgtt�����\�N�@ъ���=�Վk���!7*F�,�L�K9�^W�F����dj-�#%�l�M}��֝TrJ�)t'A��R�..�S�7$\�S��vr���֤̯��Jw-N��t�:!��W_f�c��#���1ڮ�>�ü]�>N�9ڮu�e�rֺ�9ǅ���f~ܕ�$]u���v�b1��pd���+���9�rI��V-�)����O���sQ�gL3��nIyvb��U��3v�*�J
1
�*4%`�*+�,�<���h�w�q��=m�S8���atK��,UZ.����c�?3�!��;9���噦��vۚ�9����,��_	N���|F%��|9�.}1ƹW�H���&�t�+��b�����Y�&��MQڷ�u.5F4aE�N�\������֖$��Wo�l�,E|)Z[wU��b� cl�_ϫ�~ @�S�g�()�8H�h��gs�w�iC�x��m�ƶhk(���E����~������bۓx�o�=��z�c�Qͯ��=�X�zY?���_�U� �N�V�l�h'ͷ�j
������U�ۮ[82==�E���h���~�Q�[4���pM�
KL'��(M��=�%K܌����ivm�z0��0�Ж��q<�ݣ��~���W��{��d�_	�h��5��o�ភr<�CZ�:�V��+�c��L4��L�J䏖�7%T�1�{���k��S����*&QSc�Bn���<����(�?R��.���8�QJ��q/�^�<�,U �� L������Pf��j��C�b�-�^C��1���c%G���D�/�������@�����f�Z��,��*�9K�N��cӖ/[G�9�yt�	9�y��U:ctX�b�"D�"�옥�����85-�Q5z�ݤ畲ϤV���v�+��7�.�2Dyhkq���!Ǯ�C�a���Y��t�`#z�rM/����$)2:��[�O��O����n�a[D4N��,�p�3��ӧʢ�2y��͔xi�T�+����ГQ����8�y_�q����w$b�%�\�q'*:�p���w��OQ�̈߶-�AA�X�α2������/����SYB���<�����~_�+������i��AW��eI����;��A�,����	\��DBI�}~���x�_��kA��BL���D�xc,�������1�f��vVay����S�!fq�-��"��R����d�m�G\6]|��;⿅��搊��O���~�×������y��AE���'�M{s�ڃ���YE����.�%5Ǖ�^�V��4D��f䘦ޔ6���ڪԳg�������1i2���;*�G,�"�s.�XE���u1�՞n�n��-O˟�J:�x.w�T���5
���޽[���}��)a�a��o�i@��-ьǕ毾r���&�6/��U;G�;g:��I4¯wb�//�20������bf��C*_�hɬT��Qb�L�ad>[�mK/��W�"�mO�������3�������,d8�i�mo�>#�o�?}�f澭��{5o�����U����I\�϶|�`��5�3Q��F�T<�?D��ǿ�K��CH�*����ݚ??d�>�R�V"�6�2���@�Yk�q:����l�v�z�<�`���m��_��&F|9yK�G�=z��J���ѣY�;�f�D �anS�*Ź��rg��)�������9^QF�}	f���0!A�4\-09:OOڐ&GS�gSn9B��%�̝P�H�u��ɡfR�{�T�G�/�q�a�jg�mz�M���/>j�o4&�y�y8?�㪇.�2ݠ��F�������O�L\�v���膃�g��8L[f������	2��ߎ�l_Ҝ�p �yQ�C�{�CVE.CM�E^,On��h?\��p�H@���VS����\4�!v��6�A�զ,<FPr'B��!-�h�l�����؄	�qJB�,#�8�7P��L����6�怒������<4!�;���A�M۔�"�0D�6��l}g5��H�}����	��Jӆ:it[�K^��=Օ����?��ۮa�t���W�u�3\]�y�l�g�?�9�������4�B�혡\q���M
����u��gn&�|@4���c�?ÚZ��Q8��5�� �(
Xh""-`�� �t�	�{�P�n��( %�4��KhJ�KE-!�P�,�o�����r����}�/!Yk�yf�瞕�� ]>�������G�k�����ٮW��8g�o��o�u( �������D���ƾ����Do������ml�rN?���t�Yy�c�Vw���0��e�����O�	Z��ZW���'�B%oķ�'H.Vo�o�dW=�|�=�9��TPR�A�{�_m�'��D�Ir�m.li�ξ��9������%.	K��7�>[��a��[Ch�Z�m��#�K�<���J�����&�3�Y�=s+�G���k۝K|]���/4�o���N��E�ym��?�C�D?B~SR繶����&�J��Զ�e��փ544�F7+	r��� �����G|��U���K~������
��Y�5w��^{WW׿N���#��r��%a�2R�[)<t�
Ch��h�F���)��%��Pd��ERƛ�{�D`��4;j��'���X�q�SZ�MZ��g�������Y�fm����Z餹g���?챛��g[u�d6�6S����D"VW#�xc���CCCJ�NXH�㋖?#~!�U����[�
Us��n����E��х��[�s[�:�{�1>�7F��a�kK���]��[?����|�Gq���:���1�S�k��4�v���My>���2�{>kt-��]���S�H_��������u\v���38"p�O��V�4�0��?�6�9Ԩ����F���c�,uG;�wܷ����[���<�1�dLj)�׮�L-'w;z:FM�o'�<ő�?�j�?P���n�$�lvß8]����D���/ے�ʭ�V�}��L��=��tn��_���q�n�]+�q틸Y1��$n�ŝ`�M^�Y�u[!�F��4��|��y�	��\�)��l�ժ�Μz5��q.R��}_�?b���%⽂'�-..� �cpZ�o-�S�t���r���K�W~��׻ۊD�缙}Vk8�{�řQC�3ٻ}��YVh��	 o걒;ϴ�?�i��57�YK�J��h�[���Բ\wH^��*G4�P �����!���_�ۣ~���ߔD��ZY��o��
�����P��sQ8���Y��9�/��&�L��.xݍ���� z_Ǯ�ō*�^ �s��wO��P���}�<i���ߚbD�6(kg���:᯿��]�J���i���h��m�K�m�n �e�X�&	�g��[�.>� �ڿ?@�k����I���5�-�!�3^�oEW�E��W`�$�����q�|=6��֚��F^��]�A�WU�fDHz��Z\�(�N�
�Ͻ�9�E=
A����Ӣo�Z�E�,�>]���}���E����ls�TL�*5y!k"gࠎ�U�70����C�q�~u{�S,��h������ڍp����f�E�(�n;,D�7�w{A�inE����n����Bz����(�s3�x{�+4皝��w�5/X1��ٴ;�������#����W��k"9��^@8���}��5�`+T���SD����

��SȨv��8��g�l�J��Z�(ba��%vW������t���;��p?�(���e�^�CKX5{��8ב��CV7�(�v���:Ғ7���zS+�0y�o�S���s�E�dI6�,Z ��g(P�V��P����E��"O!>(0w�ϙ�΅����������-6�w��L���n�9v�O{����m9wo��ۉ���߿�K���'�.�g�?#����F�3����g�?#��F��3�P�y����ċ�'�ط�R�6��Ijut~H���	����4M�XKN+�A�U� ����i�$a�d��I���"q�諩�7^��z�:��`��m�J{��^^a�;���R���53o��8��Z��Q�2�%���I`}n�/��ל�[��*����_����{��6�}2I~ڕ�V���oa�J���H�~�_N>�)�^�ql���������O�Jb�_�NR=Y<��Ю��k&�p ������ژ����.�pv�Q�7Y���T�&Kh�Bͷͣ�����\nU8��T�ʘ���gB�.5�V�����W��j�˯GJ�r�G����������9ݹ�V3��C��ek��7����멒ٙ�D��j�P7�V�tO��&E!CJ�@���9UW����;(3y��1�\+���c ���V3<�s�b����/-+{��kT���P�J����gB���	��y�颡�7ɐ�t�
=���l�S(aSA�Z3��mfK�o\t��Q�P�c�wU(˞�y�k��FŝC��`"ݷV�d��r�:�:�F9�*]�� T=��'i�R�j�'Z����#ز^p�
�->'�#���)��se�~���g�.r�`�w��8\+�\��������b��4�:m&<U��j���O���f�\��;����{_D*rO�c+�ttu�D;-N,��`�����D�&���&��A5t�x"�����_P��aߓN�/��O�9��7�{`��I^��R�C�^�c�W�
i|vltAS�;|�����򲺑����A��y�?�3��knetyY�G^P�a�*�<�Ȅ�E�H�q�8{��b����s���e��K�rǟ�e�����p�*�҅j������SoX\k��d��ܔgG�M��c?JB��s��<����t%w}��#���v�eC���}��i���$C{�N�5ֆ������}{�L�i�b3n>�`�!�a����1A�'Mb0..<���Bݽ?���c9�����D�K#Z�w���$Sg�o���� �rhd}]Se�k�R����<=�:-:�ޣ��3@�zT�	��k�SRo�����߯�ӽ���f�%�T����ȸB-7�$�c��aӒRR�0���2�Ҕ7J_/s�\۹�0dTIT���t�c�K�f�f��]�d�)��7��K�V������X�pr�����nX�k�K��juצ��&���<r�d۴1�����9���Q�|�ԑ�Y��d�=��E4��lջ1c*XgȨ���K���Cy^E|�r0��k�a���:�P�7|r�f�ᑁ[��N�TUi�DOEjϵ�;�D_ǜh��#�Q��7�i�l�TŐe!R�9��R���<��.��V���-�e,֙X��:,�g��(�wؖ�(�ԫ,��\�RxP�8�3���'ɞ�z9�9z���TQ�P���k��. 0u����P��Z�u��j<5m��P�?�$��6s�7�H���q���My��	��Í�m0�k��>:���o���
}]]vW<��}� P<==�Ե����'Ά]�pJ���H���'�{g�U��@+iʃd�ͺ@d�NC4�~A����G\�VT���`|JM��~1�Y�-ڌt�����45D�o�F2k��-))��g�Eo�=�n����>���A^��t��6ǰ ����K�_�m=�R]E籢l��/ь�<��EIE��xui0:p�&�Z�E]���)��f�;8��H��� 5%��5��NI��{��f8��kv�N�H.��(�� �q{{�B�����L'ozKW�f� �P�D�Pg9��
j��&�����]j�~�����uN�B����W�Z�x�����9�h�Na���9V����^�.0�Kqi���Z�����]�}ֿ%oF�ɯfXv�Q��� �X���|Î�К�0�]I�	=��h�M!9=���Y[{�I�������N�n�@����|��y�^h+��^�@���V���,�rWY�Y�%�ע�C�F�ã�
��P(Z�@����W��{/@�AC�">��I��$�>'a1��qnn����E�=�<MZ�T�P>c� HN~ ��%B�6����	�2���u�ΌP|�5���l���Jo�؟�J�`�4��R�qr���B�k�����P�VK>]�r1]�q,��������	oUE���LH_����h�~U���`%<���j������'�ʿ?]�G�ru��:,t�a����J�Gǡ�O�����DI'��⌑v��y
r����п�y
T
}�<d涹�\�E[�gh�U���2ۧ���Y3&�X?ܜ�#dh�'}怉�D��I����xG7��U#L�����5����x����-aqǰ���:p��5 ���eޓd�3c(��5���`hnd29��\*'&x��e?��t�4�-�	�j u���&!B�����H�8AQ�����_i����Ʀw���X���ZC t���9��>4j�@���oo_��w��treH @�P�������
�	�b�vV�B���n9g%�t��G^"���oD4r�����q�	�QFX�3Wo��R������ߍS��\�.��wb�GC ��)Oi�6���m��cSR��|/uo�D��r���|�@ h7td���ʆ@�����G�{�!�jTݏxE���P䌋����|4�0�uLrh�&�c�El��6$Khh(�������Ƅ`���n`�9���Ŗ��ݧ����wϭ<�9eS���ܬ�s|o|
N���(��U�%a�E;�: ���h�^R�=X���W�&k�U��酼o�������
�E������?0�zI��p�^0(�%�5���䐹o�)�����������6�0�|���Q
��Í֩�	(�g�>]�>Ud[�o��_$�!�2QGC>g�)~�L��k�@:�.;!�l��a���;��j��xM��~w��̸�Ǐ��	+˔~����d�s��D�I~��CO��ϸ��f���g,l-��I��u+$$0eߑ�AX�;KO�bn��� �	��^��CqY � ��/m4y���/H�������mr[0�_��aq�ܙ�A_�F�Eg���S���G��G�y?�л�,B�:���#`CLp"����gUg�G�}qk``@s��7�i�!��`�/��ܙ���NO���t��#��mG�B�@� ��q�ٹ����[���~K���5{h����(�^3�}�7N�����>��ty��p-�L"������d:{J�:k�6�������:��7l�ۅf��.����~B2V-d�/�S�Y/f\�Hp�D�SR�12޸q�0�+ҹ��,o��r�g�5�/H��j�`C�Y�Щ4���#����a��7�wtlݽ�:B�;�j%�$��D��*R�x<M��%��Z�4��"%�~��g5W�)]V��=-J�S��dP�E#1�PQx)��t�Oޮ�`��#�0lE�z9��i�t/�C�.��&���aP*N��=(�޸wu�;LP&�m,f��~���ZT���p!���~.�-��{fv�@��u&i����O7h0褠����� ��A���E�v�(��[_��L�"ѓ��������FA��H8�i`���F�sc�3F�B{�H$:NX�H}TD�+���C �0�	�'F����@q�]���v��u��Ӣ,��ŦbPdy�9Z)�mn���m�x�����n�S�En���������g�@D��ΠZj�DTb�)E��O�D,�<Q-� k!�C��""[0O_9φ�Z�'�o�<7`�A���r��W���ߊ��M�c��
� m�����η~�f�"�#�����Q�$��ܜ0Yt���� �$m�mI��"Q��j��%m
��zbjd�� wa���4�8J;�Y����%��`{�h���X� �hP	Pq��8��ϼaeD>vx{��J�1��>��ق��~�*�AܕsV</a��PZI!\�5$�����Ċ�ZN�\T)��~����ip���qg}����Ǧ�b��"ш�1�<�P�|<���/�[�X���W^�$m�`�2��U�#�J��B��GEu;!R"8�yLƫ��8�ķ�&)���4U|Aa�:�ͩkc���kX�#"����ƢG /�Տ�i&/�K	��ꂼ�|i-++�x6 ����t�*���	�5���JR�1�DY�v�F?+BJx+�m��w���S��e��<���'�A��N�*R��,��W�����+�Z�h��Q6� ��x-940C*��7�2��3v������;�RC�a�q`�j�@��r�f��xB:�wӻxX�R�	$[r� �B�(��`��~� :\.�et�{Z,\>�|� ���/���� ���UK�V3G@L�ڰ�p�6�������Y]�:Z;ȍ����{9F�B���~������XlzŶ��uv��W�ώ���=��U���c��������J��L�.0��f�#���~��j�j��v����3��+軗	�rߤ�_Z��6+����Z��d�Q}
�0Kx��Vn?���^�o	�M�0�#�Tw���:����s��x`lG�(������f
<�z)����6��csCW<V�4FZ�ۛ�;�+
�J�� �͸��k	)`���j�O����d��?i�CW?�f���d�d�� �Rg�h:ҥ���@��h���%2�+GAL�/��L��U(Ƶc�$�eZ�K�$�t���s���b��pl�Ed~�ǫB��y�I����XVT0WʁZZZR�����P)K�;�\<��&�QR&���Uj��/���th=�ܡe%R�@2���Vd[��h(��K�u8��\�J/Z�1��L��U _35pXC����l�0�4Bb�z�MN����hM�<��)�\6<��0����Z���i[A�*R������M�1�X�m�Ԕ�E�#aV\�ΠrS��4̥��Ol��z{g;k��t�F<$7u���{[u��@t���}�j���nA<q�5��)����EG.�Z\�<�(Z8���o)��fvܝ߁n�sn�.|&���t���\1�s?�=K���bW9U~��4gi��'5G��b���3��C�HO��Ԑ�B�!tO¯�6� �9�����γ��Whm�T�SE��τO�\������cc��K6�w �� |�д��q�D��Dd���
�Ʉ%;�Lkޡ�-1�>9�Q����x�y$"��C(�H��$�Z�,��	~�P9����p����:z���!A{nJ@5��ڈ��8oYu�E�i�u�;{�aڙ8	�����-���8Ø�s? �I���CE�-���øv=�b��OY��JD(=9ɹ8칂z7���q8�����Kx�f?����
��EW�n��s���t���t:��A�;��>�)N���N9�":��\�󙌼THq��F�K ��?<.B�>����tR�!{
��Ru��4:���8z'?X�~��Q>ц=[�J��{��9�A�n�ä^��X�k��5�ǟ�1��i�*���u�aj�7��ɨ2�҃te���v�y�L%5'����e�������,y�twPO�����w��;��?K�+;��l66<��t�uw�2K���Wx��k����:wS��
�����:��.��&5c�o��9����1�=���u��KT�̘��i��f�f-��ET���ݢ8}p�BݕE���70m�Ag]�O�0�2�gs�ƢSw>UؔxB�욦�����j4��J,�1��v��XhݬK����XqO��|�q]�nY�@Bt��������h*0Pj����~ց����
�UUs�cߜ���<gϞc�5�Nv����."��8O6��|��E��K��#S��a��}d���� �P�@�P��xL�����ɜ1��򏎿5�ml`,�92���L+b$87�bNώ���u��n���I����Y��$~�F�+Is�H,���M�zGv�N���M���O}&�" �	S��W�?�x�͞�����Y_X�>�$I��q�;Ch����,O����-���M��K7��������={�¹|�b�wQ����SB�<z�-Y���grk�8�mx;�IB�zO�4}�q��!�2�tl��eS��B�	�zLSb�cPu:��R�j'��b=�Dy��꼫��DON�v�\,��Y�iK���K�����_���@_s���~�J���G
��ز���D��Y��&to=&U3�{�1����	@�<� ��N��{�=�l�a7
w�$�3O�����t�u�y��߻0My�6@M$vOs�o�Z�JZgsnME���{/.��z� fR���0jV?����������c��C&�Sɍ�Mw���>�`��o�P�J�}��Ζ*�Ň�%�����N�V�!�(r#�s-�u,��/!�MR7���h�8:w�V� lhh ���[ �,��>d��.�\�A�,e����d(��%e�����Ч�Xy;:&�e����~��������G�f�vϧ��N�^R<���`X(ђwK&_q��һ�\�x�;����`�x
;��on�<���D�d�HL�k�;��41�(�[YBH76v3�ӱ��M2�M��s��UD#�T�T]�=]�$�e���m%�A�	<��W�{�:���Z��Nv��˟�G
����j+�?�������_�>�t��By>+�7�bz��X���{"zȯ&,���K�?�Nr�d����$�lQj��G��:>�5���}�ΔXZ�\bXh�~�p7���6�8���xa�6j��B��y�˥�1ձ�c�F����V�T�����R�.M��3�z�7zsq��ۥ��yv��2_tu�N(��^(��ޔ��q?��\��/�OjHh�7���l��5yFj{��h�@X����p������}�]��g�kYj/�����~��^�{4j(�ٱ��J�A�,��A<{�x,��W ]�/��������T���k%�vQޑ��9����E���R+.���u?C�̭ŮФ��r���`�z%q����p,��C �X;�0*%�������D�K;n�����J�C���jL��^�|j���U��L�ΑM�q.x�!#�'����b�3���.��*H�~�1����l'Zߨi�xbx��}<�o{9H;�Wr�*��2\u�|��e��0'��Nٜn�y��x��w��ٸk�0rZ���т/S��ej[ZB��>�gp	)�`�ˤ��ӱD��׳���`F�(�<�"I�_}'�?@��2Z��������/�Z��w2��\m����b�S�;o�Ƹ������%�P�R��6�"gړ{��*����/�_�?��^�sC�̽H�����cB,�[���ޏ����R��Q��A��8�:kp���8D�+���]������S�Sb�)z9s�.�>���C?����uI��-�N8����]ɳyK�͞�� ����=6;�^7)�����Q%�AG�x��I��)��U�+�(l����SY�W.��|'������%�վ[�;��ݤ��cѢ0�x(V��5X�c�榀Q���ǣƙ��îlMQ����&��xO��h���̈�(�#�Æ沼�=\�g�U2��^�a�(�Rk 诗���*�dف�'�ܳ�����X突3����}s��U̐��MoPVf��F�{�W���f�%�f��d��{fΔ�S>wZ��j�w@��X�ܱ�7�Zd�_{��Y(��RV,�?��2C�r�%x�-{	d��	}�Q/�����F�-Ϯ��ZL�^�'.���qq�T�T��H��V���TO�Қ��#���������cZ�N��aѓ�]ސ�ja��x&�Hn�=(s��}Rm����!t��_�>^�����% �4�b�!�}�N��V���_�
�jM�R��Po�������D7k�` E�{f�����dzJq��|���?֒�j��`��rn�cr���p%���W�I�6��+��7�����<�y(r����ڦL���'���T��e�{h/=���5Ra��9ob.����*{L}xDȲa��A`�Q��Qq���}8�������W�(���o%r�`}Mf�`ݻuA[5��l��\B!��p����8�L����c�l�/{ْ��J�c�":���z����!���2ǵ�w%s+Lb��ar�����g��w���Mc�&��^L�lP��j�B6[\���lQp1�D��\��u���V/�Qz���%$��IR<��v���/������a��a��F��Mqa��i_<~��0s������Jؐ=����_��&�:��p��?���� ��/�����A뉟QIz�J-�/L�����U��u��^�[~/HW�$%}gn�x��}���=��� B��ݩ�/^��G_K*Ny��o���.��>�����L_����	zh�Nx�L}ޏX����9�
�xʹ�a���
a���`,讅�N�� E��o��c�y�4���hr�;,��0��z�O���6̍DV��H\�أ����/l�����P�y x���~M⫖���0C}j�� tR�T��N���Ř@WZ�[N�ck�!���o�Ի���κZ�g��0C�荎	�����i����f�ә�Th��©A�����<�/���e���;� Iヤ�z���ز��"ts�͕0�P˻�E��`E/���aW�U���[\kQE�hш��3��
>FG+X=���v��f=��k	U�Y�c-w�=��f-�0�60�6�l%=��	b4���ߠPۧz��6=åƢ@�eDN#��4�6!��T��&�d7�;�⯌��W���.������x��54���4�y+X����8���Z��:\0lU���S�#�^*���n�����g��:�>*�D's����"��h�d2,kh���Z̑�()>������{4?*r�1��$����������_x������4]�"��Gzu"��Wm}���2��#r��<}�����s
���*}��kg��c<��&� ���c��������\�Q����$��ɓ'����1����t�z����^�������ɫ�O�N̠
�*�F���d@^@0�u��Q(�k��'D�������PnII�D�z1=��ɕ7��\Ԙ܈�g���ڮ�݄]�Bk\��7�9\�q#��������fi��Z�t��%2"Jd��4F�>����έX{��z�ѽV���.�>|�ނ����z	tr@Nfltt��7�_4^�>� {�P�-�qQc؋��m��˜��&9��J{Y�8��Tܵ�WY��Yy �u:�8��o&�� :(9�VOd�]%����J�����[%2�0�3�����l�
�ʓ�S���6����:��@�bZ��Z���wQ�ǐ���Esw��苆g��嗱�
�����
d��������?�#)�Fi]Ē�욧�NB��{�}��,�ћ7��]��y��2P�Ott�t�#&"���:� Вx�����) ����VK����j�G0q���6L�݄��gpP�s 3aQz>0ۤV� 5��{fX��y�WY��L~������	'�P|AAR�D���D���#�FFw	d$�f� Ul�\�X�R�����ojiy�}DD�m{���[lj�9�,
� Kdt����h�ĕޕ�w�z��y%w��JD�4pw$ƼkQX���!��%��,�5c�<��:��ŻC�.�d?�:�_���3��`O۬���TTT������&�8����̉�K�f�����C��@�
|y�&�2��o����O�.ԶpA5���idtF�[��66<-�A�Z�δ:����|�RU�7��^�k��,���D��B��B��Kj;�=�V
x\DӘj�	��%�	�"Xj_6�<��K������/�ײ�pts�笽:�I��K1˹�}58�\U^.�O�i�r20���U?;
�Q2���n����OI? ���=��4'��Ʋ��F���,g�ҿ��T��G���c&9H=��?4��{�؊3���t�l �[,MM�7��*6��;(���.�r�D�miQ�MN�Gh H[�͗���v��|u@�l�Nw'Z*Ox�����gkk�*$�
C>nt�����k��u��<~W�|�4��%OXӘ���Xa�"�O��[z�Mo}�)'HU��#{_h��k�h���x�����ʿ\]\䎽����q,�06���]���^��72f�*�0��20##��t��%{�]����!�f��Ճk��]��ߓ�p.U�|�{{{>�2�^�zR������b
t� �"��M���h�6��=�[Yy&Kݒ@j�(4����M����B7�����x��:|FN�Xq���J�B����?����allH9��9H$�7Fk�r��(.���9P)�C����G��h��Mc���� ,'dee}�3p+ ��?���P�eM��O���2;)�@g�`��ȏ:�(�;��E������5�^�����v+�
�ȵ�m/�N���dr;�^�F�b��g2c�B{e<�*"���� �����e�Kk�נ����0)z�9>�����E7N��W�
F_[�1�t�ׯ_�S`�_��3pBF�&QjA��e�_��J~�rA���|^g9��w�ڔ�ݛ�a�2p���y���ٟ{{}������qY�s���lgg���̕_�
��}x¨<�vD�����*	�w��ǩ�8�~u~8�7���K(�Ӿ����E+m����ZZ�;[�2�M,F��g��J�(Z�E�c���ň����t�=x���-���q��1����*�%8\?�{�7@=���$�"7S``�z�r��O��'����� s�zFp'�[��iV"����r��E�Ir�WE�"��
xP�N=}}��D$D(XZ|��@�Rjز���	G��Q����)�1�q��`>��84�V_�
+�u��m�E�R�R�2x�h� ��(o��a�t�%m��(�c\Gt�ʌr�v0�D�~?L�u�^ŰὭ����Ooa��`��-+W�Q�_x�2�<�O�^%xT��=.�~67����C3v �ƚ��ʧFQh��\,`x�r����a���f�K���j$n�� ��̬�`�%�o#7�L�Vjf�)�hM�e���������4a7W�3T����-�h���א����J#��b�׾=�����GEՌNQ��֞�(�Gh$@TA����d4}��ůI'Ckk�)����Y�#��4U�&5
#�����AT�s�vϊǶh��e�6SɃd�c����G&''�n����yj�m�(�1R&�Rq�P����E������l/�jl�"Y�y�F���3�"�1:�j�'��j�R��?j�,_��~L{}��@A*ݛ�a�%�OA��ܘ�H��i*�C[�bؕ�����l̡���nh]��	�N��zq'����"�&h3K�0����� j�Z��xJ��AJ�v�?���QX�Xj#�C$����JKK��4�p�?}R���aY� ��(�e��0���,�8,��:�b٢P��g��2�:N�����z���?rM��:u��3��P/�+J��5JJ����H��Q�2��Gqqq���9�8r��cx��%��iQ�ק�������鞆�F�z%�i�<�Qp�GQu�M�>���{�{��������"���r"��C*�'�p�x�g�N�;Uz�<����}�9�΁�m�In ���f���j�F$�-0nC��z��j<p!&󰆽ZF'��63��7}�0��
��S)=����n!Y��Z�s����
v�k��FXi���/��o-rәNq?s�@�I=�aGϷͭda�u���_� +Hu�������	w���0U:��:!z9��R-���W���Y�z/����z�7�"/�ZR�e�r�
L�=b�t�L�&�&5&��@��&t�$L��eq?�r��t���E�O@�f��_X�f��	��z�����Q�q�Q�L%�o���̀���z�\�T�����0y�*�B�������̚�L��}�9��N@FQq1��6�Y>�[Ww������{��k*�a�M1���^���t���&��-��v ��4�9A�^�9`ى�>�!8�l��h3��`=@:�an	�z@qD܃�Ku���(�>8���y�����8�Ǘ.>~~9HJE�M1�w����_����;mZ,ay�{�0rO��(%'�XM=�En`p��/+�v�$A�9|ۤS�w��H4Q�B��q�8�raL�&#�L���uĦŔ;0
����/�^�����QyB�!"���9��߇\xN��,?�M9��(�oȏ�VF�5ׇ�.|��)֡t�&^p�I~�� R�"e���pH����8˫r���������r������H���]i��7VpA�"�Ks�t������(�dV�I��|D��c*�*R(��F�6���,��P�Ȃa��I���g.>�s �R���k�"ѹ���;�v��{�����j������cSL��ʜf�\���%eێ���p���1�O��QD���*Z���%�\,�4�[�8٫󳪑7.���Z�2�C�t�V�
�)�!��j�1_��ȷy�N3�_��������LL��i���D#�R��b����i�]�#�6�"88 �	�b�<+Ao�	T�����؂�o�������>*��Rc����x���X<�(�0�uX�AQ���:�Nw@�вw=rUۈ��i
��H����V��>�\�~�RŔn1�X3�R��~�v?e��Xm�tl���i��	����/������SPDدQ6ŧatP"�'�4��x�!A�}�G	�;+&=�]Ƅ�y�\fn�}�U�C�I��Y�Y�0I=�X�*����nP������ �{��r���� �2s��Ѐz{s/]����UfM��Ԛ��0+�,���h�������`��:_F��
��> �����#���������iR����'����=є��B�LB]����%�g��ć���3Y%�
zlA����j�㏠shgM�Iq��c`~U����[�(d���W~����^@O~*�$��U�c�\�� ���!Z��ܗ��#/��K}��a�ϝ@��84��aL�ҡ֦^��"���Τ?�R۱�(���9�|Ku�@]Q�zy��ep��7�
9Hua��<����
�WɏJKŨ��T(��0�� '�:��
�Q��;�:�P���i�Ն���c(��o�Z�*3�T6�{a����$/���&���}���S�V�B$é�� ���.`p�yЈi�K,����IA����}^�pcek�t��Ɇ�4��E�@6�.@���� Ef��+82��rw|\P�/��Q���,3�hy�Q��'�˓�%87�}\O"�Z���]U�/��38�f�B�V�H��ϮK�$��[��)��qd�\͠�i�.y�V}*��=�(. O(J,4��У@��`�I�W�T�d����N�l׻��;1� ����Yy�v�S:H���bD�ѣ^`�=I��i���c�=((�E.�3�_�T�avB5��r#��H����ɎyH���v��_g��mQ_|`ݞ���8�5�q��s�msk�oH�xh/}q��[( �O-���Ϣ��By��޻�����8�Ȓ}@�y���j���w�"�7�������ܿ�}Ӝ�.�%xJU��<2���r���|����N�ow~��nOX" �7�=�����������|+���6����/!q��~��S+���H3��	��w7��j����>�JlVMS��8��}��6Ҋ�Z�m�^�Z�m�W�r<��A}�AN'���3� T4)~�NKPyRx�ǧ;8Mm�$t���#�ꫡ5a��
��{u-Yy�y%�:��8:T�Q+a�)���c�<�\���-����࿏6���8tпO?�������f<������g���f�����=����e�W� S)Y���-��l����������%�b�IA��,�G� n0`��Zٓ�	�O�ޠ��F���T�Ce�a$K�%�^������oM�?��z�Y�;��Ow�ٜ:��D�g��˟<_�P��}z(�p٦�t){�ѓ6�Õ�i��>�j����8���٨uZ��+���;����Nμ��-���o>q�����?����u�#���T������[y�N��3�X�*R�c0C�&�y��tp��	�S�}K5c�ZΥLt�3��~1as�g�4Mڦ�.�X�d�$71':=������z�#����:���B����arO V6%b�ڰ�ӿ=f��1'�&d���.�Vt�乣�%/�B�e�b�Jg�Ts����J(C�ǳ(Aul�RǬgQՂ[����[\;Ժ~��N܋֌�ĭօ��N�#��`�ׇ�G�v?u}�V�~����m��_�3�Xd:�x^�! ��f���ٯۈ|���\��i�������'c�LY�ڼ%�������t��(�co��1s�i{or �s՛���\���\ǹܞ��Ѷ���C������5�m�n��������y;��[�%�wy�g~\������1�:[�}ϯ�C�
���}W�m�d]K�r�r7G`�-[ �#T�5��r��+�T�+�$��o���E�������u�
!��3gX�����8��]ժ�`
�L`�Ė�H�R��ǋ'�oȺ����8���4�w��m*�R�RG��%89/t��40<�z�3�%f���2!��m��mH6�YN5����8��'��EC���#�ċ���.��֒�|�r����@[�Ê��#�?[�1]�+3}f�E{�X.��R*³5����
��W:�u_�3�|ТŎ�o��]&�_���}x�%ޑ����"j��G'���Nh���q�W@@z�JDS����{\��Ű���枞Q���5_���P̲&�ͺ*ʲ��W6N�����3���ɗ���;�d�[�%�T��-a�2n��0���ЯCK� ��Q���:⽃�.�f�i�]��f9��>m�)r߲�K����ҝ(Z?\�gdl<vj.?����qΈ���5�A皉D�Vg��4��c��=^XmH�bE���"ThX6��K������߮ﴟh�	|�w��u���#������D��||�k�	�z��5�{ks
��;q�Z�d�M�;J�{r5B%�|��-j3��놠&G�Qj~
7{�>v��d�H���-�%�x��gs!��-F��n����ő�����*���??D~���8���N����$���^��\!q�,=�� ����}D�Ć%R�'luO��!W=|�ԕ�e�iK�	mO�R�����N7t!�5=�O_ę{�Ǒ���뜻u�w<�����]��K�Dee�$r�K�w�s�G$�oJ.�21S�_�8�,����;�&,dt��x�N��-q���~d���s++N,H��N&�%\O1���3\m��X�n���3��D=�Wc�w��gAn��ۿ�s��r�^άyJ�~c��1�rc�ͨ|BV����r����ɺ�i�H�<G0m/0[I�-!�<F�I&Nx�fo\s�7��-?溄�)�K��}��4\�r��t4A��W�V?���H�	l�� A���m��)�3��
�6e�)%��G���u|6�����g2)J��mtZ; a�_!�"]V�:/;K5������m���An)��&21��>��Z촃{���pQ�"S��{��������Mj�HZ�����������Q�A��PPRB�i)�J����z�nIi��Q:���c���眽?�}]x)�g��b�uϲ�]��9�Y��$���v���1����7P�_���`���F7c	+�F���ʾk>���V���"��t�/y�-!�[˹�K�ġ���D�Б��cU�t�V�l�Cz}Sl��1��2��;o�"�p�|����7��{�Z�<֢乯�n��[��Ю�f0����tTğܸ���Q�5D�i�U@�\N(w��;h�
���0�@!��1�~a�B�8ϗp���B%�ت�5<M��5���]��h�D�(Z�`�Ax��P��zck��g��Ci�G�ই��Q �:���?�&�䓶<!�P�����Vb�F!�����x667W'ˠ�ȾH������7��X�ma�^-�#zP����2�Z�lޓ��lbMA�!n�oi#{3����f��6k�D?��_f	`}%�c	L��~sr�lx=P�F���NJ��u|��?�{�W��3���VҽfN-����=;CW*3��^���a+yw�:�\��̹��i��H���6>�!�6Èچ죛��e��M+�7�\�\D��V#DWb2�f>7�����C�#��~؁��p����(�.����SlF�
'F�`^������v�Y�3G�:��m�^��S����Ϩa�y}�0����Lk����k;�`�I����{��&%A��An���:w��^�c6&�\�"(���l֜�|w�l�����!�B<MRP�/�DK<nZa��vx6j�"�������,���v�t�J޹?��۽����@����2b�ҽ[����s1���'s?�+��5d��P�+�Wp�)8J���<�;�����e��xE~����@�&&�M>��B�:l,FU���v�w��}��M>�pd-�����.3#��ejb\�H��Yo/�RY��`�M��t�+��8\u�7h:�+�sh�r�_�1���-��e��j[����A.iB�q`�
}�X��f=Q���Lm���S�p�?���du��/�/:%���-q;�:��ݞM�lV`��T�]�k��Ih��®!�k<e��̷�t��U�[ڸ�È��9�a\�u�#A�݄Z�v	ͧu=A�Z=w~���$�i�H��@* �ӯ:/�~��O���!�?a���w-����69�u��J;>�0�8)�u����Vϟ��(I@o��8S����Ч�&�������3;%��q��^}0φ��f��]�$T��{�o���9/jj��k�())D���_��0� d���۫��p�1�kep�a�D�qZu3�G��и��h3oiE�~_���a�N��
E��������?�[����"q�N҃-�Ӄ����u��:��L��z�s��]U�6�>`�-�@7j:���w
��{>��C9��IHZ�h>�N~I�>�)���ֹ����{dx��*)�:��4A�=�l��"r�4����O��w^��i^)����h�{{�#$Z(�!�5qIkE݉���(.X�����#�*�H�]�堙�hҦi�\ۊ��2(�c��-�<�<�m��GE��҄;c�OBׅo��{�A�c�F���|����E�h'�ɬ�H�5ٙ���_&�)B�Q��j!]Kb��н^('��
��}��& z��o�v�Y�c����R#�ת�̨��F��Bd��{������g����w+�}��*�4���+�b楏��A������*��*�n�f��DRX�Û7oV@�|%�����R./�Vk�v5�=w�
��e�3����^F!"O+��ج�����yN �z���#}��ÓvZ�I�n'�<��T����z �:�Co�r�
R�mD˩&0���IH~��S�����Oޠ6w�re�E��x�D�q����^Z���h�u�8 �Q��[�B'l��F�$(�K����OS#��DV���b�#��!��c��<#|��%�g�c��/wL����(��u]B��q+��_5��Et���t;�,Qz3���t�غ�w��:��ֈ)�K_N2w�I�j�o�)qCg�u�2"�,[m� ���'�7�`��:{53���a��Wm�������f{�҈Av<�i�4	�b��mippG�� �[AF��\���jI��y� ����.��&4�(��ݨ�n�@>8��}��)z��p\���#�k�r������0�Ƴ�-�J�{蘙���m³ȱ˕���$+q�����[�2�i��]�ZO��-l��­���0��wKzԡv���D�����4m��D��V�]�w���)�?Ox����H��y�AY�B�n�#��Ɣ�SJ\O�5������;�������c��c�/�D��(�������8�/�=�c����8&�F̭bn«$^�����͕<f��;N[����I����������{{��dA_I��Г���Zb�=�ݐ-����K�U&G�A��%� ~�D\m�/��,����_��߱���<f�_*جK��~��VR��y	�.B^���&i&v��#W���#N�9ی��MlX��g�13��'��ʬmYxm�yIT��ʢ�a��eǴ�����q�8�~�sLݑ?���B��6~��d^\��;�>D�L�����Kq��@�#"��=溴�����w��:��na�X���)�]+��z�a�j:��]��Q���L��-�%s<�j�a[̓?.>��ò�_i�ѫ����FP��+�+Mn���"��l:�"@���H��q�su��JKBQ3�Ej�A"��OՄc�C�ĝNs���P�,��0	����������lbĠ��0A�V�T7 %�M�%�pK�]��2��z%��!.���������|�g܎��i[��R�~�u�gU>D8y[�C塗WS $�%X+[ѻ� zݮ��(}��s0����Vt�ʡ���q|Y=��������Ev���Ν�#��mF�Wq�� ��quM�M��t{���>V�y̻�ٳ������o��E_Eb����W�ם��0d�ꔒC���i��xeT',�J+��_U>fI���T�����c��%koE��o�aj�-%_q1�8�+�>�f�j�Z��V���0�z�7�sAB�� {���޸��q�ֵ�>�CE��E���o0a,ikɌh`���U�m�3���V�'�M8Z��6�_렏�Г�?Z//��*j�:�z�������i�Ԣ��Q� *��H��|]\'5���#z61����C����	��K����5�¡Ew�y�����Ԋ����=��]��։��e��7a����=��;�7����|��=6E��'��f��ry����Q������1zo��/��a���9���4	(S�ZοJ�K��_�2rom���*|S����?_\�'�{����"Ӵ��'{!P#���h��8W�G�k�r�zMe�>{�_�!���XZ%����.vb%�mb�e�����K�-��,zuJ��+����a�E�jڡ�%�����d����a���%�P�ŨaY7�wdߋVB�F��N��q����+�� ������mѴJXNu�#�U"��tӎf��>������`7V�yq\v��\����'��3sֲ/a���bx�D�A~���Fv��~��Qat$����ɓ8t��p�<�k~e��߯V���;����%�B)��^s=YE^��&���Q\�����9�A�,1R[�{o�l�0|��gK{�����ی�g�T���_`7�sssu��~�*k���1����<�6��9��2=�C����>����f�!�R=es�������2��-�����ׄ�\����������D�=���)���Y���N��Oג�~�����2����9�9�(+.�B�!�V�=Ά[�'m�X2�n� �ռ�EI2,;�Ƿup,z��F��H�*�����ltgR__Oi��ڷy�=�>c�vٚ�ڳ�n�c3uQ�[���^�]Y�����X ���Z��������-��e�bc_t�����k����a�yX(G��XOUhw���/��ǫ��Lu�U��b7�������U.˟֞�}�]a�.�I�7�🟬��p�8��Ǜ�X:�}a"p�e;(v�naj��t�"��w�kH8�pq�?��������krrK��$?X��=�8���6
7f�Q�Z3���
��0A����'�J��ݝZ�U��=倪X�<~��Q!��.���v�j(�H��m��.���߿)ݼWz�?ji&'ӄ����_�����|TW�/�D�8:�]��
8sMȗr�_�'��Z����¼��j[A�p��N����6�D�k��>C$>�mBG����Zr"�^�}�����i���4M̀��+	���Vq==��{߶0�P��������ү߿!��S�ȼ*�\%|�����|����	=c1p_p�ND&�56>�c��}<?oP�[u||��]nbѲ�R9uu
�����,~v��@.��N�������O>/}���N���|�A�_c��Jo�&6A���Ȩʂ(�0 ��DST���&)�/����`z9yy��tX�T4���o`�����/8��Dh�A�nB��cՏÖ����x���*\���B�>!5HR[SC�{j�/�4�k����M������E	BDJ�?�-t̶���@#�mi�=mi짯���4�G
Khw5b��2Yr`��\�JH�^K_�� �P�+z�����ǭ��efe1Y�Y4��A�=,���?���t����9�M��	�t\	�"b��>��ro���a~1��W�on��*keU((.�QS#
Z�]g ���T�W5�Ret�Nh�u�o��ʓ�V���s�������D�ůr�
�2��gVt���9���|��9Xh<n>����*bU�RP�S�q��!�[�D��C����U(���U÷����Ͻ�ELv��z���{��p`����MMt�׬��Z�qj_8к��AX�N���C�A�f+�
b�}�J�n�^�)�SdGގ�����5x�����nf^�F?��i��\R���6���_��ӊȸh���+��·�_���x�A�H&�hV����n�(�/l�ud�)ſ?�� Ȣc��Sj��j��zzz�[����uLѼ��]��)���nd�k<S�ۓ�߻7�3�&���
�VmX6>�-�J�Y��C��ׯξ��M	�����w������zG�Z͋hv~�Pggp���
�{����)*m�9�πp>��� ���Ѿ�׹������K�%�p92���on�L���D�K}�C*����ecÇa.a���ޙ�F���.?�Y\�Y����ĝ����UR�zʗ��d��>8��׻�g�R�-ΒX��l��OW� x몝�U�v~F'a���(p5�*tl�d�x����y��+�ߨ��N"��M��֠���FJd�d�>cv6�VUdnKZ�q�{�X	�LѽB����'�:�����Գ�����S���m,9���C ��f 8�7��0�o�\>���-������ǌ�\�B���a�{%a�۾�a��Թ� �4ek�V]D*�7?LLN>O�^$��s���=�i�u��sJ�����ۖ�7f�J��{�Q��(0�-��n<2��i(eyJ�|q#��.�xy:�Uf����$;�y���O�����m��s�.Ð��y��>���JVcz�3b'����>+fudz8��xD�<:�?��D�@���F�b�����:��s��ݰ�A�+\�f4r�D����������s��%8���s��-Yn>�]��L��E�{�yL�2��GbM����瑃��h�G�~GI�?�  \�ݐM��eVN�

|�0��z@AA����g�(�DQ���9������cc�F�Z�Ω�)NK�)�E@E/ha�
��k��#��?�D_B.g�O��Ij��WwOJ��@�|7d��S���}U���Q7tt�����C��T�A�*�ۋ��}a��:�2	�i4�v+��Տx�V�T�3�#e�	�εi�����q�ړ���z�����\��nS`�v�㠤�D�������Ų�-x�w��N�lA�������|K�������<��;����W5���`��}�������s�qf2eeecGGҴ�4a�B`�o<X	 9�(<�����X�un��l�e�gs��wu��>��J5�����\%��w�J����`���T�MhM������w�gff���ni�MOw��N���rȃ�������]�n�U �K4��<HT�=��#���(����ebb���:_�G!#��n���X�)=#cg�4M�$�?��w��ڄ�����x�ܷ���	��cvV7.��G��K��F��r��-,����]�XYY���RV���tc��0�K{u��������-B�A�ju���x�3쩲���GY�����d�]��:|���sWCv��S�TѮ�+ dzzyc�&x٣�7�*��YӺW�I���h\t�&%� R~�}6���B/c�}� `�����4���?E�54zc�r^�����j����l�:D��S�� �pg�m�Ǐc�=:���y���O%�NT��SS��X�ˁ�RRQ�j�m�}��|�3����Zٛ��Hy������"|4F� 5I��֦-�Ť�6M�6p����>��6� �B<Bm�b	��k�U������P�x(���L\\(���n��2�+a�F���
�mi�۳��]J	7����as����Jh�5UyPhZޘV�?�= @8�G��3�yJ����ذYD~�:����>��2�|�V����5�;~m��z=z�jQ�܋��6_�!d��~�c�:::�؞����y���\;�ֆ�UfM.m�p2��T�I�����w���&������3����b�ى�����R��y��v8�>^�+��۶$bG8-�w&(���2���:��;� Z|�>}��'��pp��
`�%--و�E�'%QS>~����&���M���! ߳~+,<�2�+�K��4��@VR�h�s���_���'b��|� ��Ϡ`�����|�z���hd*)�����aC� ���mJDӊ�===+�g���[&.��OU%ߎs{d�)�}���-������8�����?lz�%��D�A�`��`�XT���O���{�BAQQ�L��j������mfFۤ��3�p����w��B��fL�|�9���
?���K$h�H���x�eT�b�� F�FEE�B���<e`�sw�`H�8/�a�z���m���5|�ry�JLKϰ��nq�\�o�a�+�4�7sqvj�����w����FB@ �?1��!6NG��C@W����+�|�����N��"��e�A�������=F*c]�o]sZ�4���-b�1��4��,@Yz�v+��׌�����ү	~��L7�x-F���2�䦨� ����� Vf��t8_��Y88p�����1�t�8���"Ъ�m�em`��ڹ�x������Ռu9h�UCم/ꍘ��Ϊ[h���V���3��mYs ����t�Q[�����N	��H!Y�wM���U�+͚ &`��3�^ž5�y�!�!��lC��Y��בm���V+C%)��*��ͩ��������l��n< �^	Y	���~�|d�^_�VYE��.��R��\�B��B�Þ���?�l�<�Zn��\�E�@Zt?��6��
{��~��to,7NM�~
ȳj (�x�0OOO�"{o[A������H�M��
���m׭������W~�[]3�<q^���ZDD�h�;�/�F)v>�.����h��"�SB��@�@�$i�\�u����qg��k>>rX�ĺSVa!����r5�]�=Nv������s���\��R��%E���� �D֖ȫwrD�e��J���nB����E�TN�w���5��Q?�|���z�/��������P*�7BF,�A�u�,��wS�o�_@�t���E ZZ_Omy?������4p�zUx����fǆ�m��%#���6f>9�B2=|X�Y�MKn\ ����P�����Ƽ�==r�FT���~�*l�l������`h/�/_�6~�w5σgي���WM$���.}����H�b}����mR����m�,��E��f�6X���|��[��k�	W370=����(���`�tX���3@Հ~=�NII�0��� ʤ��ɝ���v���R���}�=a5�$O[�NՖ4�����؛�+l&_�j�:5!O���OGgf����B��Ê�lj'g�/�%�/ĪG��� �D�:�(�U h�dǌ�)�ix��{��C��ͩ`'�p8l�
2�"��BK �T(�|����*3{b���"3���?ggg�|�I}����䫊����u�4#�)�/~"3�48b@��.�NJ�7f8�k���ܶ�
#昱�b��u�h4�r�^^��I?�gSӎX��=uu���tm��i��/v�Ps_NU��o�Ke��S�|�6�4&˄&nmoWl��,��=���kB��8c��1���6�6�y��2��~�_��̏	��x�+*j��\�L���¢'�B���-��w7���8��v���
w#<�
YNЄ.3��f\�K]	P<�7���ϑ⁴u��4�5��^of�,29�=���T�}55_R�=��av �F� D�w�����8кh��`����؉��5�eX)��ͬ0v(;��#�����c�C��-��{�xR
�H���k(|Fnjc�w��;������Ņۼۮ�ʛdmtMKIn\�(���;��6�)l��Z��L[��zl�x����� 1:v_ |�]3-hY��){Dw�Sϸ�<�큚���t��M���lKE������5Y�+��v�uTb��I.^���0�_��bWztjҀq���N,Ֆ�PFmڂ��֡� ��3`26���k���R��?�Jn&==x����L��b����.�ݲ^#ԤAA�VG��N��\
�+itcc��\m?�&66�+����������N�b~ʕ>�j�L��@Vs�
�S��WDTT�ɡ�Vw�2�}!�6��T$n��b9��?�7{ ɀ�}?Q�
�$�*������LE �����?���G]���$�'�yҖ���WQS#k9M;l�w{T�#��ˋFZZ:�����P�$��C]�Q:��
�`yy|����(#����s�s��}�(�/���0(���LF�Ջ���b�h�+.�eok�]\�]}��c�DF��Ur����L����"�����+.&$��z��H<�Pa�}G��gb"�b�%�f��#2�=�"�d|�3��aκ��U�:|Ř�j�h"�c���Ғ���'ZH���y�˅���+4��X�z�_=�X:v�:���׿|�O�q����&�����F�A_�PR.a�&j�(��A����.?��&���[;�-�ڹ/�*B��:� ����%�.���EX,�l����]惏xƘW����s/1��Qŭ��� �G�sE��m�BZ���>xD�ś� u6������|������.\���s�l�9/���T�����c�o=~hʂ�yj���V��U�jݪ���d@�4˛�t�y��qqqaMmĠo�"��Е�g為�vfCg�}��=0A�1CF0Թ�٨�=��E�C77��Y�2�p9.����ُ::OA��^���a�z�R�(�B������s�Z<�\\�?l��'�}���}P�ψ��;��ի�%�m�Q���b�������+m<h��h04v�5qW"�Mt3#d��k�����VQ���C�C���p��r!���!O3��p���0]�v^�q���ݳJ��`�ط	�r��^��6.�����.�}tw�4�Y��}��̆7�?�5ޥ���!�aC�mhH��df��φ{���{׹�#�����ռ��-~�L�I�_��B�l��R�]�����t�@� }~�Uv�� )a����oM�j�P���s.�����^@�b�f^�I��͞�{��T�ik�i��`�؅cC#*0���KUӛ��Z�hVԮ���������b��7x�݃AZ{8��uˁ��C .����y���ye�烒�O���f�wx���r;>#�G2p(ej�\__'�%i;Tu���{�������(*���*�-������"�Y�H�������� ;bs����6\�W{�0��L�Os���b%�'f5�}��gu�����Lll�p;/��L������_�z��	U�j��֟�hˤBY��v���zVr��%�}n|8��Ҩ�>H�L�g����n�X���+��)_��S~�����߂���!6�^�q�+�Plz1T�	���
��Y~��H�QSS�cj���\���#��� ?�-|_��{&6��`Á<��"�뛺M�<���b�)͋�u�����\~�N�f:���a�임��Ą)9�?�nt?��D�˨�	jJ�6Ͽ�RH\\�rK$�=!v�n0YS�{�0�Jj�O�"&���0�~���ӯ�l�CL)[a�g�����,�p5�ә��^^��E� ����Ιæ$�@=c묘'�4ika����T�o�̌������[#@�]5�s��$�!�=M���fV����T���Q�ئ�W�ܹ���狰eض�H�-��w^)��D6ꇈΗq?	���ee1-o(yz��^BIb����#�_�2��T:��Ԫ;��K��zɕ�;uxH�'��:rNUij�����"�e\���wf�Ó���y��k<8�ɬ������p�!_��St;n��UG�����Ӈ���A,&)q�Ra��b�l�2�!�Y�#`��/��⾸�r�'��3�x�r�����H��)- īE��ؙ��<����LO�ۡ�2KJ��s���0ޟ�>^��B�1/�$p]��A1��n��M�(~lHu���?z�s���p9�eJ�3�t�`��n<� Q$访$�m~
`���)))�W{?珇D�����}/�W����|C�C.����VYY٫K	��� bz���~J9[Q���R�GmMMǶKO$��\K#6�y��W���+����Ҩ�>���ڔR��S����wUz��=PK�D`ve%9 ,�3�%��R���tL}����;�sp�spp@����V�>��M�G�����UY�` ۨih�f���JCC��١KV�J��f����@��5,~i\sJ��i����O�Wq��/�P"9`��pq�������� �+�W�-_;;�o#�g<���/g�4Tç�_�
�*��;."^�J�߱�����AZ2�=����WoOK�1K�k�/���o[��>�g�ڟ��ي}g>]��}��$��ud�>^��ު��p�M?*;��Y�|�軐���<�� �1F��B�џ�ѳ�²����r���G� ]��*HM]x5KM�h�ZM��mᥲ


Ⱥ�
2�ī�F��ws>"	�ˤ��h�ܣ!�}���V2'rwE�����]w��vyJw�.�k���I%�Ǒ,�aB�!�
�?彼�,d�2�~@�]��1�;d.�gO`��D�I��ĕ�4�L�,9՗>���9����\�N�&��h=�<> ��\����ޗ*4��MB����>Ϥ��XZzfa�m��C>V��+uM��!&��������
�����y��A�o�~������A,@r���KJJ���t9�2+�tbƒ\����%�pq'�"��^1�~PUe!_.�Xq]8�� ��� �>5e�;U���Y����̈́�TҌ;8��!؁s�G"jٳ�`,���"�'#"��B4��;n����Q!��{}d�7�_3�;a��&��3+�����ʈS{N�hϒu���d������H4�:;�<�3�g�ѯ�Sn9>t�,r�Ӌ�}!V}l~���x[ś�w�,�!KWǫR�VUZ1Q��ײ�`C�����?H��*�;
xF.�P��[R��Հ��fMKKc�E$�iሄ�5m�ޙMDD�F���� 
 u|d\BBNe%�����N����m�i��;��]ۈ��g ��[V6|&��]	����$�>,W@���z �-�M���Hi����o�2�Ű*dloo���$�}�����Ҍ�4=��E�҇,�m�}�@�w���s4��_	Y��&ؓ��:|�g#���M����}#�u*1�rP3�t#�n{}$KZ
BsQ��������$��u�ܤ�r�O�oA�go�R�ckZ�8�ଚ Pd��&ओ�����rm�k	qت[���;V�q���u�����7ge��-q�6������'bo�K�}6��1�ED���^�Ukv\O_?�r�
b��C�O&�
�S�W�dC3�(�{{yMצs��y�0 ��-4����(g��E�D�*&6-1���d����H<�67 pfm�W�._��d?��h2�=1#m0]İ)��֦�tu�[:���� 7mr�w�9��﬈�����怆�).��OL|���y�j�|��?6b�.	�-s'�-Y<<��	�մ_�Ud^��mE����i�#�RWg1���y��l_�حlh?��F�$'cϊl�FC�Q��]�b���Ғ�L�(l2bW�&�Q���=lb�X�_��`o7&-*J���rPnٯ��s}R�hr{�'i�SUs�[5M�|����(��.��6kg��;P�gd^�`�Qat��c�H�Vxr����(��N�r�����)��3��-V����
;T)�{#追bf������n9�!+�jZ�\�B�y;���22A��'�{�|�*��������6QTr"��]H=@���(0�����6U3n����?ޗ#߁Iw4��V �#�P� ����O}y�ԍs
��w덄4�ձ�[�'���DJ��i*~}��{a�b�z��T�jq�0k����ݡ�QI�{��V���kf���R?���M�%���1�xx*�Qg?߂������܍��~hb��� �5R�c˪��VF*��|��#��Nf�@|FFFy��"]��~�({��sz]��>��?دbٟ{�<��"6���')�P����K�����EE$AQp��P�x�����\�d�&��v�!��g�m_=A��F/]�7�����W#e~�9�ҽ�����[�J1A[z�� �������T���f���I�ܗ��j��k�Z$`!K����]
7q�ۜ�?��Ԥ7��_Eyߠ�ߍ�/4��	i�4��"Nym��u��W�d7����$7��m�l@�B��~��?Q��ؼ�g�վ�e�V�׷o�"]�܆BJ�ǰ�W����4<���'��o	o����q#�8���55��������fϻ'���j@MSn|R���K�[���&��hh��f�f���զ���4��LՊh_
.����w?o�9�w �#�j��&�Sx�1�BKw;������f:�w2�=mi�Z�޷���q��B_uG�I�T���=� �Ζ�������Ξ��``���l�-ED-Q�~�%;H����
aJ��4d�	Rp��^,�un#e0�Ve�E��z�A�x�q�z**��߿����a߾�p�r`o�n~�U��<?�7�[,(x��_���Zq����F�I��Or?+t~�����u�|l��'��O#�F9~'kg��C,�ꋼ<��0��_/�g��T���rmE�]qKGdI}/E�ϧ���H��G������Pm�kk�"�����kO�ߔ��
c�`0�
ȟ"�0�ͨ�961���hV_}.�$������^�c����C,��� 2����[������5�M���6�%��%N��$%q%��$��� �qܛ~�%h�$��iq�TVV��Ɉp�$�����Jr%C[�*���Ύ����oe��{�ju#s�s�bSs��.�c��A�B�e��~��.�UCSs�l{<�l��:ӚR��X�ԩ� ��H�k^��c"�����[^��7�N��+=0�OÓ�I�f;qkn`�K_��,+���u��󊉅mo[�b�j �����f� ��B��N�}���� ��q�kc�bbcc3[Z�o����30sS����
��)��K��U��g�c~兓9��o25\:��������tp�2����**)��?~M�-q�9�b�:��5�hat��
�P����9�SSe<=��m-�?��)>��Ȉ���e�t����ذ�c�{��>;�g����.ѯQ�E����yZ�f��]g�
B|��9H��L��o�π�&C����bb��߃��������6�R6r>77Ǥ0s�F�&\J�R���$6���Z����\)���d�aC��ӑ�P҇(���7s����T
0!��4%s'`5<�~����/��/�v)�3/�����=?�ۛ�Q��dm�74�`���㹎_C�J�h_�WW\�������wdj�EAv7��!}Q{�����'Y�{Z�����{��_��JN^>�8=���:�8���/��vIdp`l�$>�!^z�ط���D�6��Lo��3?�@���������ׁ�����X�K'dI���!z@��vAF]w�#abk�\u'K	����^vkMX6{>Lȕ�x2;c�	F�Qō\��]�f4�*S���cjz��b��kɖ�C������ϼ�o����� 
 -1c����B�0� �yW;��wJIp�@@^��J&!3Ǟ�0{��������]}ơ���64���kD^�^/���d�fߟ�-T��x����Kw�1=�'b:�;��弼�i�.�>�l�/K+�����-md�2����ڱ��M�p�p��^d�!���T�SPP�2EmR�|6�,�p˳��Z��������d�E;�k�u��1b�!v{�ʷsJ2. �VvώR����V�>��5$�4��e�FY�׍o*�� ..0��>yw�f�dr6�DZH�DҬl ���re�7�*^�W�P��᱆Z6�� %�J��-� $���;�K���:�����������iy�\�V������{]����-$�֋U%�b�aU�q�B��UU�A$��]2T223Xg���8Zr8BhڮfI���HQAO�s�8�YS�^P���<��Ԑ��=���6´T>�X��w ��Yϭ|��:E����|��YV��3 � ��5l`O�`�k1�����@��g���h�~M"�� }_%�n<ܸ��C���+p ���+�S�{K%���*4�466V�{�}y�n��\I	��|����Q��(��X��+�����������A��D��n~^�����2��ǀ���O�W������^]��=���2�Hp!~�6Wm�p�I�}�<~���s�S/o�c�	�=��f�KS��Դ.�����%���5&���&�6�hѬY����?�+���#㚝+��qd�n�'��< �#���d�e{M�2/�Kj���ဦ�-�9�q����7���55᪝7�ebuq���{���P�ұ�{rrB[ 4�
���w5;��="���e��ݹ�ɰ�!��e����=7��� ;P��/dk �i[[c�6�Т�.��w�Dtz�A
������C�����)�B�,QNNOV�*k<�t���eQ��DO#���*���;�Z-f%e�i�%������9Q�g�ٞ ��6aߕ���Ybkt?���v�������Rw��>��jQ�%n9Y�{t����7���M�YM����6՞H!��`�^��n�/:�w��J=��kr�K���|�~aj*�(�ۃ�<�EE��*�!l�+]k��Y�Տ����C�K-�vZ���uu�Z�s>�����ۗ���K��lO8-���Մ��jX�4Q��c�hAw�:%�+dV5s��f
D�����F��fΎ=?W��sÍ�T�q����g�z_5ha;��K��>N�p+"xǄs�b�Ҿ[� #]Yxӭqtt�	(T����jj�ep��Y��JNiM�NoWm�6��n�i��XY���봭{=��8�w��s-D�O7����I�"x����^4�VM]��L`����R�444�o�R�; I��+;}S�JN�P��	��?���.(,�<�.x�'�S���N�A�0�S�+��T���A�`6�m奻��o��pՁ��&���ٿ�q<�7�O(�)���.Ѫ��JQ��B����S]�mlLC[�A��3$��(�6�Mx���ӛ�����O��A}��y��ރ��wP�,[ܯOb��j���h�E\6���Rp٦ �n�=��=_��6�tv柝�S32�x�F咊sV��S;u�.!�5��S* �A��v������Qԕ��mq�K���6y(�df��Top��-U���UI[�3�u�9jaaa�vv�����rÐ���\\��������CdI��N�7��k��on��3���;³�����7���]|C�����2��P�,U����_�����:���͵h�֖��G\� �ֻ��i�EEX9��3������TT�䮬���w𝔹++I��_dd�, ��Ȅ]��t�@�>b}��iVE���Ń�Σk�c����۷���W@�X98`�e�C�c��gH��P�����j�l��ν���'E�loo���'��D�J^^��_�2��TYii<=}���y;�+�B4�Wi7�k���@0U��b�Ҡ�ᯝ�g�������S�6N0�J��o �r�TE�m���=��殑�e���zݏ�wS�Pk�G�n)����D�a�����-��꾷a��A�E��SB�FR⡻;�K@@:�S�FZ��C��w���oƑqn<�9k�uŎu*�.��+�����I]�YXX���7�s���qt����$������E'd�ۯ6'�+d����u���E���?s3|�Nslg�Ư���,o����{dWk��k�Lu���7��555�Y��Q��(�P�xtB�Ռ�9�������
�(�S�{X��>O���?��(���86<�]��*`9���G��Y���1(�}k���=�;�ׯwo���`@��g��������QW1������ug?C	q��*A*�����Z�ۻ�mfo_���̀�R9�,���Zvi�W��H��;���zr�P����CG E��=����Ǫ���qlt�
%u��V���ޣ��̋X#vK�\e�s��Ж�fT�%����T!�m���\<��N^�;���0ҭS�R4����,,-��U�m�ڟ���ř�e�̷������属-��PR���c>]Y]��6T�lVM*����՜s�ʊP3�Hg (����8�b�ҥt��%u7,D�V{%#����sk���jP��ݫ�Z���ߜt%k�Y>ZukIqu�S�-.EiY��d333��<1�mlk#��V��P�s�PqFD4����`�A��t��9=`�^��SV�Z]m���d|������@�!���ڛ3�ۧ��؍�[[Tbbb��@��~A����3d���-6�[?N���gpX��L���MK#6��+�.���ɉ�9�+J��ۛC?8�_-�\�޴�%)-�S�����cc������j�m�,Z���C��`�7��Lv(.x��FpQ4L�(�n'gg��{���r���8
�`*>>�9C��/gj�:|fQQQ�7{3e���g#i8�e��|�����U�p��]�X��~A�Ni�a�%��#l����f��;>6�ɡG��7\�ʾ��p�8Tc�j����ݨ�����O|&��.:U�}��Hu���ܷ��lnY��Q3i��ɠ���!Q���Ekǐ�z�ذ`
K�W*�j׍}7�B�����{�/��r�`�W�3����,?yN��8^����'�]����=��ֆ֫�R�֮}V�""�>�������Ņy��lᒽ��k�/X@2Ì�Oh�MT�8Y��Ʊ`&��0��]���v�S�D�J7*ӿUZ�U������"k�Xސ�lSE��ܪ�/��R�y���RSX<n��05?k`��v�r�P_��F*�D^**,Ċ�J�Ɯ;��{�5����W�;��_#|+߁�K�~��l����+0&EMO�s	��U~�ӑ�g��T[��eϬ˗�^y{��^�k���S��n�@RM��UP��-3@��:�L�z���rtu�A�R$j�- &	�s*���Ɋ��&п��88@nǩ���8n���}B�n�9�?//�ܕ���h�����o��ϡ��!3��Î�]���艌�oܑbA���c����"�Z8
��+)aRŇ飯�>�q���o�C����k9�I/&m�/-��o��'���~m^�;��}󗂔�)�#S� g�+
�ȵ�="�*RzA���^����JF�i0�B�m�C���������8ϖ%Bs�dQ��ؔ��(u�|Iy��OO�,�s���|���E2$]]��ي�V� ���姞+!��r�ͽ��7J�'/�;`+�����2�EMH�uU+��o��T��<B��m:R-������*.���K>־4Q������N���	II�@vT-��Ny�#�m��O�g��558	�Y(�8��3権�8��u �ѧ�:�#]��v��AGgy�Y�500@������А<�A���i�̸�aǷ��9�U�CujYhU�sn��C-r}��תj �BBB���x�!`���B1|֌�W�_�ް�M���z�Z�f�&�z"��k�矼UU��!��`p72�w1e��+E<�j��# ��Ny�B���+�Y�Q�]~@�������� L	���y��2�;Ǧ�CD��g#��ӨV.�L ��*%5�C{Z1��CUE���� )���V�߆5gD��tTF�RMaiupO��L�8�*�Ə�(�Bݴ,Q&���(ny�1|ձ\N����.��Y��A),=-�z-�Į�E�pPl,���jY[[<}���¼ee#���
\�_�z���\:P���`
��r}jVV�J���{ը�]=��CA�I��M��ll���?��	�@�P[]����16~~شM�#I��А:��o��,)44�r�KWp��痵}� ���w>@w�U��d��_�}rr2J����;?�V�KQ�7�����h��kRz�	y�IҔ�)����0:rK�>�O��:�UQ�>pkɉ�]?^�%���%r�\ԋW�9���Z�w�0����*�@������8u��c"���H-�c�����I�)��bb����xl���\G�B�e��v:+�2�!B�''X(�Up_�nf���R|+��QP@��4������� ��vɼc��rkq�;��b}�b���?�~�{�Ԅ���R�!%I_3w����o�%ɶ��/45G�,�c�M��D&�,:&�s�읩)<P�&&&�h�/A����i8����g���������VH ��k��B:�1 �����������IN��k�E5���c�H��q۷����4�V��VU���ч�����q@H���T��y�������q�5��-��cN/`w�=��7!t�|s�4����=�L��t�o�����%{,����n����\`>@w9f:\Tȅ®��<�|>����O�rJ/��Wk�j�������s�7�JJJ_�^������yK���	�[�����w7$��1,-Բ]��j�ͤ�����rZZHD��\,-���:�����deb��\�?Ivh��� ʄ��hH�36��S]��$�e?ػ�i��|��7yY�Ka����t���;Z3�k�q݂��k���Ύ��WH@;^�1�{~�4��"�Y���Y.��@Bf��[��������O��� �F}:�F��W���$1��W/nօf��	a�L���8�,_�����Z��~]����Ibh�^��}q5�S�P|�{_�K����ll}d�K�P�~�[�XR� �"�T�)�#���IZ_�G��a))a�]��Z?JY�s�/1��S�D�����#���T /(��ZgY;�Z �w+����K���u[��_׼�5�ꩬ��tx�������o�l�/Wƿ%��Uʓ�Sh�
��OJJʓ���4��O:��0 ����	�GN� �EPl�ywV�ɳ$�u��k��M?r��Dd�+�����se�fQ�~��:#�[��M~<h���I���>����R5��~|a!����i�q��Kc�&Q ��#*\��:�(s�^��M�E�������}\�f�š��DR � -"��r��ޙ��6�9�'�Z���!��r��ɠJ�uޏ#�!n^޼ϟ��]���D!.E�����P���;���A���i�R�B[\Y�&+$lx��n�tS:���g��i39��V�;�����+X��۷���l��򟪻}�Ԥ��^S)}���6K��s%gZ"��\���� �ﴁ<�%�*�"�"E$��~e<��x&�o�����N`�CXj�߰��;>A�+�ҵ���+k�ɜ�>)���6�t�9Kf��Z���9vh�tP\ZZ8C����W���ϣ߮^N�ec^mz>�W�ۓ#t{֕w���^^�<<4͵��%�����)�G�=ɀ���g7j��K��Y	�~���չ����J�:�=`j0����a���۸�̈"�L
�3��
Nxx�@��Ij�=O�766�YG���	��(�"`��&|jJ���I�,	��,8DEc��*�23��Q
������p�������~��Z���r坴��:��s��N��KL�F�3m������]!��.���"��'��[%��*t����(.MSm����g�XC&��#�^�	DT��#��v�Cy��@� �n�Iސѯ,5�I�-���� L�KL\1�!���/�� �x��%}A	�	��������M]�|��Jz�,�=��ߵ�-˱����ZZ@���Κ��tQr�Qq�7��fWy%Q�+W�ik%����e���}qس_��0h�z�J)�Y�DcՎk��{���Yf��u���wՄKvV	��'C�DD���0�dGu��޾3����\��{~���o��D�4%��|�(���[��DP�|y���q|�g�UD�b淛�T��|�-	0�7i��9W �_:}:u~���g���Do��Ѽ/_��y"�I��E�(�`�~ m�����TTU����S�Y�\L�	���x�T��4�U�)!��B&�ֱ�WT�Y%A�#L������o�`�^�mf���f�9�y'�o�8�����!��������JEpC?}N����o6(���!����	3��vd��N�O�����EQ��4�[U<К���<4�7$��4Xj����֪��|2=-P�h̙(42��'J��q:;:v8���s��sW���&�ۙ|�!�;�����F�{Y��B\��K��}�'�2��5S�ߵ���&��ЩbyyT�
Pl����jSd�s����@�xq//]q����q��ɨsIձ�R�3�Ur4D�*���&��4�x�!~׽�;���KK������\ �񤢢���.t�r4�W��b�;r�w�CI))���ؠ��t8�+O>��f�T�F������䚫c�j�D���TM�q�A<�Z�w�>r�2NA����|�Q�3P �걆0�T!�`z��о�9`f:idU��9U�Kף�	�q3*|I���I���n�F����xC�/���7Y}C�/�R�j������v�5x6ǲ���s%���Q@<��I�J|Ս��#����'�g >��66�4������7i2O�Zae7.n�Sĵ�SR�[P�yc&Cɽ��[A��PJ%W ߽�0���bM�]C�CP0D$P捂��R�s�P�`ww7!9y�[{4�����g��GҕI�Ʒ}��UUW��Ҽ��A���|�Ǻ~Xh9ݩ�<��;&�	��/��z�/<�56�&��M�5����Z&^ӒٵW�]9���8���:���l"�e��F#�+'0�u$.�j�A��o.0��$>lQf8�����43~��g�� �sѣl�XsflX�챢�8����rl�we��c D{�������j����͗\3�Ӕ�(#����������VS�u*���8S �yq����hQ�r�
 b_��"�����8C�K�%{�J������X�����+nv��*�r"@Ct<\(H�h4�۪�3�f����Q�i>�݈����>��ʳ���逸��Oן�7w(;�?������10jV>�-���[�X"'%}?�R�Bۈ��~��H�/��{���Ó�!B5/"n[[P7���	� )��ޥ����qG��/<:�4ssJ\dx\�֌��ܝ[�ve��?���r+,Q8�O�L~�����-�Sg3礥���?&&�r'ڪH��,P�H_�����.^_Ù���R����Rz[�4������м�a�A�l��<�ܮ��^��ܕ���[��=0@�v$###rl�[�:z�<��%q�e�ܚ�*������QB�UCA��٤_ثl��]]XHk�Ҧ#��Cpv�le\�l�kׅ����䡼������z��OS_����_S�k�&`Thl5����+���m���Dsh�69o㲤�F�ӳN*�k��JCC3��"�Ðe�i�N�w��,�����4h��j�V6iқ����=���P�Y�R^>*o�C�A�+EE�i���]��qJ<12/�5�d^�2��E�/q��qzܗZZ�Bs=��g�r��a�S�%�$t&�dd�WVↇ� h�����2
>,��������k7̴����(~�
jOn˫�m:=�B��swu�H��Iނ�J��Gqd8^~@����,A�����ڍp�=Wx�С_5���	pB�Ȉ4p[���[�s�	���_��\Y����m�������(�v� &�[tKN�=���]C��U	r�UKl���o)�8z��������B4�eЩ��6��F3T����	 �n�~wN#�%w��}��g=W9���s)8C-�sM��t��n =L'��[`Ʊ�i�"�#onn6��&��G*�!~:�]`<99���]�m��}\4ĉ�Ũ�[��mEs��\Cdz-n�A���4
�DcNH�f̣;%��P�lT��c1����5��D�z�;��i��~�[�&222����ɾT��AcMAժԓpt<�ӊܞOM�1W�l'i3P�5�8�8
HZ6�¸��}+�FI�h��&J<N'�(|��u9F(��S";�r��!o8e*l���BzҪ������x�Z&�f'���2�-l�zk��+��25�t>��Szzz�����@�����Sd�����ܓ���I�����W�@��n˝
%Xl�.}�"s���p��'���e�����,�C����H*N.��Ag4|-: w"�Q̰��#�R �4�47�|Y
����E+3�����BЬ�637׽~L�۾`c��Q�Y��H4t���Bĺ�:B
�㤈��2��=��Xw��SSp��3�Ҷ�g�E5}�k�&:�����e%%�?[��t'Ё��nVۯ�^��.lHc��T13vrv~Vj���.p�&th3�aԱ��$�Edu"b������ޝ$	\�n_l4���V���v�z�|�8�X��=�4b�N��ZN�� �@=�P�콅���U ���krss��cqo66L������N��8MmiV���g+d��F>Գ��w����eJ]ޛ);����ck�|�f��������ff�C~��t��m�d��Z�^RES,M�}�GGq��N����/Q�?��x���*��Y1Ǩ|����b��Bn�fC}���X\�n����f����46�Bz���u���5��u�U������5�^k�� ��D�kvi��X����>#�\�x�T��a��IS�~D�V+�W����闢�"y����tt��;DT�x�ޞ7%��X9�+e[��%<�M<-ԏ����`FqY�߯��a+++܊u���їz�ys�/b4���T޾��"`c�e}�uǧV6S�'1.$i浴�T�:"��G���� ˁo��f��F���Z��F��>�&���E�n !�� $�p��p�5��*����7���s9R2��֗BP �ց!��a���j��YLi^/�.c�:>J�.Hل����W~~����	1�
�=I6�q�;|�+��ᯜ�c��>�>�{�RR�Q�gM�ީQ!�C���gTe%�������֎3�e���  u�]�0��얊�o^~�x���_�T�5�+�g
¾M�_�~��q��Od��UhF�Y��	�˔m�fJBI��}�ۈ��� XZar@�8�E�xR�SW���=����u&����ju�ww�rJ�N-D�[L�CJJطo�)y��#� ;^��W� eSM�oo?�V 9���,U�@@�N��-��^��g%I�?p{�� "���?�%7�-��6�b@�5 ��A �.sa��8Զ*�Ȅ������5�E����<�$|�x�P#]5b�����jM�/T8~�����9���}xx(C�+����)��6���XyE�ZadA	[9�e�'�7s�Ʉ�R�I_,�Cʇ��2jj�y�J3�}Ts'�,-w���4$�R����	�d�ۗ�W�����`?0�.X����J�{(��W�GZTdd���	�씐�R�'�A�r���{~.Ãega :G�����[EQf�V�|=���P���6��Bf||�����MSI�����e/_�������&m�di����7.��n��TԚ\D��i$@�D<2i����h,9r�"�ꦖ��t!��x�#��s33 Uh�`rj���T�i��}���Ԓ5.��6o�����H:�R���@�?�G>H�W��}q�|��w��w���t���y���|xV���9�I��,- �*'���ݎ',W*�?O� .�Di������@Mv9����7�%����laa�EA,UAZ���Hc�9"F#<8(��d�	mل�㻵pǈ�������T��Nm�����@$��j$@��!��>b����55�[%����Xq�bk)�Э�gԸ�#N�s��,���f$ԒS3Ԟ.}�7��k>__N$����U�貁�.�ׅ�b�Ap��.g�B�|w勋�?��ϾD
��HWz1��,�{vh(�l��ۦ\Y0f��ݐJe[�������� ����/!�V�Rg&������I� l��ի�߀�	�8a"�p�iJQ�3���&�f}�9V�)+G}!�����#����������:ؑ϶P�Qۍ)�F=H<iy���(�mF Dm�/�Ό��`
9wLf�+��c����Tjp�};��e�-P.-��[���)�r��T�͝�}�����I�j�-��u���k�����K���D����{�eUU�:���%@s�=[qH�����k�}}�T�m��iQWS�� =O����o55��E /���7uhR�
��� �,g�8����8�_������,�k	m2Ҵ�KY�Z8��	�2"��'�%fw�)x����_��V����W����^it\"�+���zB���������п���0r���J��C�*�Ғ�@3IQJ����@פ�_���O�j��b&D�)� �y�"�qŃ�jRb�י����RFBy�܄⃨b5I�p��������104�C�����������C��i�hUG����qP�5�"iq?
1o)��N�$�,�����ll��%�hfq��Ue �Cf��pFӒ#<<|�q�Ă<�����$Y�=�<-&�����5�Q������\�}O��e�7`n���#t�XR&#���T��Á���J�����C�ex5�����ZZd%�-��gZ�!'''4��#������95{�lN�9�a��٭f'�/L�-7~��[������FHV��|�������f2�܅m"�d�&=�MSV���`\����͗u%h��^q\�����دξ�װ�(y���[_�9����{��1�I���`�a;;�McsK''l��W�kX7 `�r�V➞>WA��)�If<��>�iii����2�4U�e��H��1��-צ��Wu^^�<�1<���1�	b��۬O��6�l�}�>OX��X�x���/�^>��<#�E����^�����꽻��{_�3�H^�Yn ,�6~�g^����sU)>�%�J

�3�GGG}3eZ*����`���(�o�U���������Ē{q���<���j�f��F�M����i�Ҳ2�eU����]\$S#�6�/�L�||HA�V�d�C�K��i�q��m�Ad��^ѹf�tEIsy��4I��	Í����+�_QCt�I�>:��!ꫛ�7�rs㵖��(3�sku�z�[ww�%;�7�� �O|_��9�թ8�×�����a�d�-ll�]Ї*2�U��>��HS��%I�UF.R����w�4u!.���!�?J�-~�C'��K�gaa�O�����߿���T@*ּ����0k����rRt8!�\v�x�3��<�_�]�@~��V_MMM�(+�����|���t65�.{��-#cԤ��ν+��(��|:�j3_+���@8$܊x��)n�:ʦ���2 ��233�}}}�e#׷�ԧO~���R3윔��#Fy�4�GU04`��NMo�� ��;��'�i6�|d:�����r���$�_X�A�)�4*��8Runl�܆e�����*&G鋣����C����0�S�ʪ�U�	�9���K����r��O}^M�j�U
*�RÍO[q�/H6��
]�
*e���iR�k���r+�:p�tL�j����}iI�gˠ�̬V��W+u2����f�m��{k��X<(ka�-&����-'V�������puU�J++5]�y�04�n�V9Z[3��n�$�=	F�B��z��S}�	�~2u����W7�h�H`�e: %ۯ�����3!�Q"��P��F�NS兾�,0~��=ɇ^��}�4�i����kt����`�*�� �B3m+��KAA!~1P&�"�v�Q�Eߧ��7��ܿX	*�E���F��|=a�gF�ګk��}K�Q���ԇX���y�+gzܮ\�0��6�<�f"�eV��m>�O�{�MN`��,�
rs%&p�i����#��A��������XD2����Tk4�gX�b�~LI*�e���5[�� �qu�G^Mu�50q^8Yg0"��5�[��
�����-<��v�Y'�:�����0O[k,�6��j�Nu)*�'���N*ޞ����8WUֽn�/�����(�r��mͼ��sh��i�4<�g�`�h�{r�?��Tز���؛�U�oUT�L�6��Ĉ3ss��E�U����������o�tX�q��n/{�����9j������
\$���S����/����9�}7��K��96vi�3��v���/�Lԇp{,[ˈ�ƌ#�á��h�ρ�˲��� MԭQ��(�V[QƮ��&߶?������A3Q�'^�+����1���7'��1N�o��ճ�+��2����4Y�AV0��m;� O[����SJL_�u�32HA���L�?�o=���D�^�&�F�Yo�����d�IYWO���/ ��y�󍎟�N��;a2�kX�� ϶t��������Z��x��X%4�7_s���%]c��/0]m#�kL1�%)^�����gez��b!&gH��nCK���!�ԏ��je��
#z 5���#G�&,� �׳��G/��/|y�Tp��n��k��s$#6���$���<�.�bl���,����k6M�S�/��-����^���eƜ�o���	�^�WI�w=1)q�a��XݕG��qS;ϕ\���Qebd��m]�aƗM� �-�iw��������<�B�@�S�P�-?;����T��U\^i�\�̸�G��++��+U�K����h�iL�r���p�-Z[[�;f�-���"�wL����(ur�4�Z?^�Y8�Z`�N�3�O�}�LϽZh��_���<.�M��Z�Q����D��ܭ"�)�z��(���t�3�+�XZZ&$'�V�֑-�|�;y�O|y�������U/`l[�Ưe9���%��c�܉*'� ����G�Q��t���XD�:�I���o�����v��R*���ؗ�X�i��%vvV]�z��R�s���U$��������i��-��W�����h�@� =���k�V#���
 j�┅RSeUm(����韈�tOA���������T��U�Dk����WRΪ�G��*6v�����lT� ɳ���y����M�e�D(��*T�hd���Ţ~/Y{���t�<zh/�H�`~�21	ɚSU�'��)�JP@(����3%JJI�s?�19*_ι�T�n/i��2�%Sނ63�@��(M�����S���3�tM[k�Y��D����q8A����I��P[`�`��H���XY5ˉ\���؁���)� ~���n���2Jt�˲���S�{�Ղ��D��b�|9�5�o�oZ8�p�����d��o`��ؑ��W���G��� ӗe4��Z�F�9X	ӈh)�ˑ��FB���лIQ*^{Bc�P�4��s?m��i��k4S�@����Z��T���b�:�.f�m�g�Oګ��]F����y���Kp3����P�|b�!BCP2��X���g+
~�ω��>5o&=���Y��I�+��zC[������p��O���oX������]PP�E>>9�zF���t����~��Z\>��5��cm��ZUH���?�4\&������v:*�Rn����k�Q���w΄�)���,�F���𐽚<b
���l���Q#�đ��U�ԃ��Ы���]Ϳ�7��ybU�|q���7��p*����e7����J��dx��D�4��חvA N����ݥ?��o�����e�K��w���t��pQyP
�璘7�	�,�R;�,���d(NZ���"О}�/T�P�?�3H���f�u9]9��X�Ntrv68��7k�X�m#�lY!\��\-#�F��O�J�W�U��=��v�A�B�;s�.̀�7ͩ��ޞ���t��<f3���z|�8:���B�����x� �_S2%F����Y/��r�C�����P�_��뫜5l&ggǕ�3��1�����obbbaa�t~s�qشmD?Ԥ�c�"
Wm�2p��L�^�×�l���7���*M^��(��s�-F	,��E3����g�V�NN8lm�T-���w��(�ӻ���/[(���)D�1�����T�1߭��D�f���yC���
܇`��d�Q[��5?~1���"ֹA�jm���T�YYB�-�l�/��-{m]�'�}�VV(����í�k�~�12'M�A��0
�h��Bk�}���~~8N�Z����⇋3[���X�n{�����b)C�K�1���j6��yS�Fu�4l30���*$<�f<n~7�_�#L��;u@���H�9��*�~:��Ň�����%b�������f�5,�5-OO�F�Hy���>�x�'��u�q��P�߉�MA5������H5���r��_�cޙ5�F 
1O�t��� ������j;wT!�v[n`{Z{ҵ�,}%%E�ݧO����m~-��۷1�.��w�9t�9��*YNurv�K����jV�k��X��T�U%c��j �p{�z�#ҩ����Ήm�r�)|Rx҃��p{��~���݊��ʒ����ů*��}�N/��׺�N(Ј��HHE����;[����i����Ɗ4Cc1��"�O2r�{䝐邑�F�D}܂ہ���#�,���n��BBn~4x���e��e\]]��=�h7z�����V;5D�4/�<yO�?��:�'��T6� �2�NNn<�W�&5Qu�5��D�Eg2�P�F+gfvV&�f�������x:��
�onf�"(��5&
l���ꖂ�׆���ߪ�)(���Kʩ�w��/���,��݉3�W��CT5W���gy��7�\�>��EFg
8#�eH�f/�L��}�Ŕ�?y�E���f/��ۧ���<锲�o|�ch��L� J�^�2rq��7.6:��OZ��T�������c���ۓ�����On�zƪ8-sG���_Q��x����Y�?c��K@����Ωoh	ѪGƺ$Jq�8�%�z��$��'��WP@GDD�j���u�������]�M?Qg����|�0(6���>��l�� zQ/�~TQ
X�5�~�=�����(�v�5�� Zm�L�In�3#���Ů_����8K�0F��5���Q�䬦7�Sރ��i����oŉ��F<��q�*�:�Ö�vkџ��jm)m2���hT�~����`�o�~��k�fRT���w��^�:�<��C�L�f��!��E�~>4OI�Ɩ⓵��d�x-c2���zrs��w�-���{<�ق���(,d� ׉������x1�o��q�$멈��?d�P�퇆�|~�.v�P�����Y���`~Qۍy���$�zF̈���Ϧ��
l��u*ZZ@��f���N*����a<���(�Z��o������4��,�X��c�����i���Ӧ���z��+Ր�Оw�o ����B�h��H���2}�g��W��4F2W��3<<��R	#����e����v�Ҹ|H#bǿ����&��BGrV*1)��[Q�)����k%��
4D�KQ(F~�b�n���߼W�7���t��?�0b_�	/gYiދ]th�z�L@���e�s�>�Qj�DI�¢p�l�I��CE`������2�T&� �������g������9�0ho+r�u�Y���l��.�ަ�>0�r܏�m��j����M��^2�LI�:��T��U6в1�5U2|0}�v�SA�s���vFT�Q@�ڇ�	`$�C�����'����w�Yf���A�ЪRZlF��J����ᚡx��d�E�Qns��D\�U}�Ѳ�<?[�i���@o^��g	�����8"������)�c��w<8��&��{F2O]_���4�x�G�̉�x��<�n��_C^��X�k��6��*�k���6]�����̞ɚ�u���?�U
+��2Z��L��_:���U�G�|���vr�)2�c�XC��Q���Ι��߳߿����|�K���_k��"K��l}�|����qn�s~$I��{�����Xr��G>�d�%n2���,����4�<|���)����J��c<�ZFn�Z*��p1S����Z��%�1�GtDɥ=x4��(ꠓ���'I�M��Mӭy׼~;M�d���>�_.eL�q�E��|q_��m=����!Kl�D�L_�1:0W#7�A����sz�x�L��������X �+�8�Ͱ��;�#Ńlgk�sw��@L8g:P�aJD����dΣ��*���dC��}��=lg1f	�׆�-��A�	�������b�ʸZ�W��#=i���N��V�g/)/GC@@��Iw��G�8�>� V�>>�w���%�U$V�ݬb���k{V�h2���%�码�y��F;q� ���X�[&b����}�F�}��m�"�T�E�-�'�qq�iԫ������jd%�m2�	+�1�g�@�5�:Hͯq�{�7Q��hh�n�����8e ��~�����"���ԞjvV���
�Pk��F�I 	���vI���9|��y~�!쉓�L��v0���nT��.�mn
Cv��*!"A��ك��Nt�cY"Q��a�ጭ�#�{��^�	1l*���1׳��v��Up��ܡ��]5-{�]4���1.zII��޼Y�-��<����I~'���J<C�p�Jhz�
��`.���ҳ�Vd�ӟZ)&�98kv�q~h�G�N1��157��E�X�K�P�N����N�j#�����#0_�g^4��P#��iqͲ�/�����"mr�01��s%����"`���_��V�Q�m��5G��K������F+ѝ�X���vv2JJ���狳у;j�-�o��[0Up�NG���(s�|���-�C+##�G�����4�������Y�f�`h�&�a�ͤtl������y##<�)�s�l[�#>25�s�ۼ��D2�����
(�#�6���b�՘a�
(*��jgv4d��8����A�q�ܲ���������?.���\e�I�:zVV__ߥ�J��#���\�r� |�H�k,x`k.W�1�x9~,.'f��o�=�?f�Lˇ��w�L6����2^�}������s~|< ���u�g12%��i�X�u�;.��w�J�l!���+U� e�����q�\�h��ŏ[[����>�t��"K��D�_*-eX+s���]�d��ϙ`�3�5�:՛����c�ǘ�����k�q��,�=֡�����!y����%&r��P`Da�'L�L��-�v	�TS������8����|�AB+�*)�lI��w=��'>���@�ro*:��~����)���);�8/��)�n�Z�iK`r8->ԋ`]Y9�:��+���=���r���-���*�ꥼ�ֲ�Ԕ'��sz���8����2"N	�`�n|VV���M��!%�7g*��{�5���� ���9,��R�P��z���7���Y8������> acӈeAǦuc������V�YPص��O��n_L�mBg9�����TW�5f'��,��ᡑ���-�d��������1C�����c��[��rƮZWhƮ�`�蒝����)���D�juT���"�ņ�SdXh�\�%[�vOm�c���d_�-6���,;��h.��H�i��Hۀ�KMM���Sh%6(��̬ӆ��Ɛ�B��"���ݼ�JV���9�>o��C���Zڷ�u\#�+Lӕ��׀-:~���eՄp�ֺ��w����	&HW�G�pc��ũT/*
ʟM6"h���HRE��ʹ"��\���T�����#����\;Dѫ�_�7G)u��P��0�"5n�4�� �`������@o؍�,R�s��u���f1���A�,l�袈W'��]��Y�?b���,��j��)��c��1#��҃�HN.|������oB\�~w��q��ᆮ���$��Ze��=�L�unYD�*���e +��]�O<�e֯�dBj����>}
�y�i�pf�m�۽}������><�\�MdMhQ�z� �@�b�,�(�� �ê�%��s999)��D@;U.��13�lr��jLU���IH�;��>+փ���H$ħU���B�V[S�*�0�Q�^�ĒvڜLF��I�O��X�C��gg�	Ѻv]����d>c3&Ev��K �$|��C+�2p����^�v��?�g�o�L���<)<a��S��x���9llU�I$w5
��Ɍ?��u��Q����*>��J�������Y�8��*d��Ԫ��7ݠ��5��L���
M��6��{-/l��W"@��00�aa&�����貿�N����ϳ�~��&��b�f�����:}/�	Ϊ�7��5IO�I���xrgh�kc�:�=���N�$�/eha�����-�`�!�!�f�kD�0f5��i��J�7y�!%S�[�����J<-�7�_��W��F���)���5�:�.�A����NX|t!C�f��<a��OU��p?m嚯�2I����N$
)�i�&=�����m"�{>��^֕��'�5��#h�nU ��'8�)J{���s5W�ø���c������*z��o�3L�8���_;�����1�0���#��(>��\!0^��*)�V}�z����<��8&����Dl�
�VU!�f�tܸj�r�Q��#}
�`0��joCg�>����?䞜�̙���B�U$p�f�'%'�MT���G1�X��p�9�+���81�k# ��;�J���������]( , xcs���{�7�҈G8O���t+�y�XJ�#JK!;::Z|m�g{�73��!uO#��9Ȳ�Y#G��q�cfJ_���S��Z9i����N<����6�V�y�z��R����tW�{xl,�7�����kﻃ�j�6PA%�  �H��T� A	2� ���� ��J	CP��� q�9H@��4����}U��ڿ��ݭ}�nz���O��<�i��n��EO��P�,��R�|.�3�S�b5�@3��� ��-BvD,�8XPQ�Q���i5��S+k6��/�BUBpa�Ao(h�?b��_4��z}���E�w))�{�����sa�m��(�շ׀��q7��2A$�#���-+�At�w���-n2�1;>:����:�a��фk)8����!?wߑ�Cِ�b0ȹ\q&��yp�����d<c)ߗ�-w�{�J��Y,��<�ڪ:"D�Jޣ�OCK�qs"�pfNK�pesݜ�{�O���]�)JO����������%���WW����:��r��`Ik�����D��`�y��Q4u�[6�b�o�͝��s�2B���@�Q�z� w��s:O��t*�ݣ�L���祥���%�¶w�o�*o�������)2|��2��NL�Q�Me-X<�w^�mXXzb&-�9�N�N�#�*���Zr2[�I�dM��/ݥ�*%�>'i����dg��OK��!>�غ\���Z��kr������/���Cm�ӈ�Ly�����,|�z��!J
���w?>�}�i��eh�*y`�		k�]!�����4N{5j?���䐿<@b*�:E���BZԏ�w�4�����E/o�E@��Q����K��Kg����u���d�[?�+a�A�U�O%/���ϫȃ�E���Z%9@��o�h�l]�WJ�-����ܳ��*�yF�73�t_8�)�I+I�%���P���#˞���m#����\��_�
C�Q4���X��Ո�6�6? �@`q2S�a0l/�����O�I������H99��r���R�/\����c��w)�\��()-�6+y���
��/5ן���h�X�ӻrN���}R��Vh��T o��b�gdsgx>=��YK���dhhx�`������x��ƫ�v�f����mji�]�iV��`��U��	�PǤ��X����-[����Yl�/$�I�f��O�z�0�j佐���;����fVm�����T��8��뺻���c�K����Y�?O�3S���Y=�ɸ@��o9Q�u��4�dY[^�	��
�u��g�6��l=��\���\{#&�u�N/�/d`�}[T����9�[�%}�O^p�U�f����/Fg���r?~�,�|�M�3�S�~��*X��y�`��P�O넾{t�/�&ԡ��zzz�V������ܒ�7�����Z�շ���������7�|�۲��}���BU����[�A���y����*wIM�nر�4�ꈼEZWݶ�n		q^������}�M,mr�M�},�v"�js�!{+g����M��g����IZ���ƍ��8��"4M1��{����a11�ܔ�ܧ��M�b94�D.4�T%���r�,%��;r���AJ����o�q����Zr��6��&��A�����'����Z7��Np��g/)vc�\��O�ϑklGM����\9wGUUu��H@h�?�)�/�����x��7��T�&64c�^�F�q��P#V-V���gm*Ն�A8��B�l�S���n��������M���]���A��i 0"
8�]PMif]�ҾBe�GGN�'՝v�r�*E���6t�ϯ�ύ���9b���O�)E1��X���zs�p?{��t�lD[^�E�$)7�\�q�3��Xt�c�s�߈!](lcZ�b(nIk3E�^^���XY���ά������m�x�\v����9 �nB�L�D�6�p}�����WX�k��e���Q�y.Z������M�m[K�!G�X2R�UHS�Poxi�~���k3�/���55T�q�;����R��]�9[�4�9����*u�aT}�C�f�ze��]���@pp�bK�/�M�N�
���A�p�	ǩQW���?���0����8j.3�v����%L�Н
�&l�}��0Té�0^�0��KnW�6'>����'b$<����I���v7��.^��g\4����=�4�v�r�/�h�����
U���p�Iֱ�EqA��������RR���x|d���<3MU����n��𫦼�w�JdI��*oU�ĳׯ贋9S|j�3x�e��/0�D��=���fBz��p������h9'?����!	�ڒ'��H�����l���p ��#S��Y�s0:+Yj`rVI�|sCC��w�9杴�!k!Kfh���|�W��Ӈ����YS�q8���'c�Ԯ��D���ҟ��-ќބ��O��;��=_�6���wu\?<��'=���rG��ؼ)��O����N�1�嵗�0�*�e�,�L�v��(��|iY���년��./����&�2 �������!�[��/ڙ����b��Ue���h��b��$Qj�7���w�;�0.��#�Z�����+�h��7���?�9R��^_�h�A^�����p�1?�ZUU�<�r�������(�s��Yg�#ŉdWV�j�p��8b����3LY+~���p��3%L'/P�!�Dݫg��Y�Q�Wu88j=��
�B/���H ��A�B��J�!UC��0��34�$����������o�|����xx9ꚜ�A���@�O?��b�J%���nJp��������>B��%@,��+�]}��b��Z� ��Kz�wXA�:@� �Y�T��Cg?�ߩ�8]�pbz�Ò�;�_<F}�S��Ǩ���d����N�J���Uv��LM�{�z��ēf��~9�j�R+��|M��߾��ֶ�%��2ņ�䯟Rd0�ki���v��di1sf��݂?�\Y�Ys$��L��3�,�2�ï�d����G_v\ϟ	����gG��e_��r@;Rg�-�O�i�8�C	���������N5�팭W�����h��3����^�e�
!t��KnOU�����ξ�k;鵵�qO���{��V-��烊t�F�hAYP���837dJ[��S����W�#�=79����=*�UK�V�'$�y��*'�f��>�o�����(�d�������e���N�v��i��1������A��j �m�����Z�MV�
���}N���}����m�S�F����|i{YYY|��[^�S?N.��ә�$�9�,�?��s�4�qȒzx���4ɚ���A�ӳ�x2<y��wБ���[s(j��5���s��L�	j3>
Z�00iܘn6ÿ[�z��-�w��Ƕ�W�����C�x��)����j_���?�Ójc��7�%�	_��cC�?W��t}(|C~��"%>*"<|������緖e�Mןy��-r�l��5����v�e�q/�t�z��y�B���Y�ǩǪ�����j�x[�|��>��ܘ������/K��x�W�[�����b�H��,��_�d�ۗ�e�iD� ��킩�"�4k�[JA�wgx�����'�����ꄩTmLMa��o��'֚�(7@|(>j�~�]�����	 )ݶ�+�TW�ƅr��z��`�|ɨ�~t�Tο	�����۳����ljjj�7i�L=V�m�nd�cbB�L�����U/����_��Js�1�g�0���[��1����u"?Ǘ.��7�&C^O5�b�.:o�d��$[���"��iLLB�	���z�	��7~�w�����8�$0	U�zg�@��X_�Ǭ��T�*~�/�![�-���uz���E��n6XMr��Ϭ,��)����zC�|�"�oXr*Ϡh��Ή�ͽp�8�F�{'zztj�3�]~��θԂ��+�#�ON�}��������F���N���s~�x�{	ZMC;�w�[x#4�tI��M5uuk���� Pk�DNg���Д��P|�.�mc����f5���S��O��i�l�X+}(�|�"9�詩6$���|u����W�Y_��ؗǫ���9��$��"�O������_�$���Ă��N��O(w�*�]2��>T�'g�z����©�̀�+�Κ�~$HN�XM��MwMr�y�f�]W_��KJ�;����;e�+���wutz�y~��כ��>;/�arr2���ҘWT�vd�V�n���J?��M�����eS��Z��v�Bϯ\
�z�|�wB��ڹ�+��ܱ��;� ʭiA�y��Y�|a\�P�qhh'��T�忬��ʹ:�`Ɯ���l�� �jL�M?� kP��g�?5<�@3��sc~��|�̫!��5O�Z�̀Ȃ
ϊ�}��
S�cs�����dZ�@����;6F]�m����u\Z8�&��P���(*����Oi3�~�
W������rSsT��th����Ubݕ__}����K���R_���� +k��@�6�O ���3N�{ܧ�C̰�̑ryWY�<�ϝ`6��������@�o��j5�9��ԊV�J��&u�Nhk�&�_�/^@�5pq�%��3* �}|H�Y��&G���0;���W�㇤,�6}���n���1{�$�,#��B��o��U��禃�`_��|R�ʥ_ ��b�z�(bbcc�
������$ ��r��#�|��QPi_�R;�`�X9�Wv&�8���Q�ߢT?�$�%�1��>)r��e�UzEI���O55�}����oL�\�HG�<@'S��q�k�8T�Z]��q�0�R��UQq�ߓ�A�E�̂9?y��o�_���&�ȸ{���>�y��LU�Ж�HH��+�~>��
4��z��4���7 e����ʅq|�ˠ&	*�5<���y;sZ��\f����:�ӗK)ھ����b|�?ύ�4� �ڦ��7u㿢>7�������
��x.hJ�L^�"/..���$Oi3~�ڪ
���zxxX�QY���eIg���q!I�	K��%�"�)�t�U�AjЫ����ݳ����Q��	��ł���\�/:�t�T�ղ����o�Q��;�'&"�ހ��=iii0��Q֫ka�����m�ݫJ�b�^��+�/�6����[�B���q^�(# 9����u����`h��m�-�[Ё�P�,BI��G�=EE�?��f�,��.������?�n		Y�����%�[��
�Zu���J�֌iZ=3���kkz�+�M�g��Z�+�V����t�����p=/��nK��&m8���j���Ů��"u�u9���3>��-(��Zg�ߚ,��֪�����'���d������D����;wdd9���^�}�+�h<��.��������K�J�j��:��Pkq&s 
�Z[[鎪�7$9��t�]G\�~ۆ�E����kb�w�I�n���@��1��U؇��i'v�8a�����~;�Y
O_���P��x�~:h����"j=q�������_T4"��uVm��Nܻ���g�'}�@�.�[�P���1?��ʁ���Vqe�cB���>�b����(1�*���[����t�"�¨����nk��AW��?Ǘ>�y�K��w'�j��F�DR"�
��3�8r[ZR����ow�L9�&����6G'�ă�:�>raǇ�����r�3v�z�]�INW+(��N���	����?��:>���@*��df=�u�pHf�x��'@
�� :w�'o#�J\���>}�kkkˠ^�z���h�ׯ��P�M␉���ZJ3�o��O8����Bzx�����Gyo��r}��2�|z#CL�����X,�SM�]�k׸���1��CKO��J�J�i壽�c�5�1��Ǐ�-#cJҘ��Qu�3ͩ Y�轻>ߡ�mO�N��l�BG%]om�F$g���Ԣ�,O�w�K���ߐ߆i�Dt���:ZH-�l�&�G���Z����z��>/ �@o� ��WMߘf��+��Ϸx������!����jo��.1<����|8���������������F����?�ܿ��rʷ��9>������.���`�c����K7U��Z�ݜ�_p7�:Y�x�XO�$\�-��M��jA<n`:��/ak��yΞ=��a�{!�Q\R����X��s���h1h4z/�x7ꀄ=��'-����:��Jv�C}�{�<B��G���
��!!�x՜�g�"�=S�'�L��/�d-����8d�fƽ&p��{�5�ۣ	h��bꀃx�ׯ�@���rq����I𬶖��N�[_���ǭ�:zzzWW�7���''��;Mt6s�')L�I�K����MTG��W�4�3-���pmm����cv�m׃�m�q�)����Ԩ❍T�u�OuH�M+��z �<'��%	�&�7<�̮�
��r�iE�����㠣f���'	Z4��b|$�Ǉk�@���1>�e";QC"�t��a�k}��^Q�Μ]b��|ŧ��Δ�>�;�ܴ���5W�fw��2���K�5︮�RJ�;p�l����V��ks��}U�'�z���8�x�Ǳ�\ve)�N�h[q���OV%���:����L�i0߅��]���544\fg?�r�U��G�t��M��Z�&NV�qK	�P�(� �BKS���Q ��o#?�\��U�m*+J�u���c��%p�K��K�92'�晰���(�
d@�
U��k�j��;��45��F4=����&���2�;8 ST?�:�<Wx�."" �+�����J����`���Byi8��Gy�}��}���*�*�7��*��̬*v�y��4jb�LZ�����ph��9���ŕK�� �����<.Зz_Q�rz���꽃�.7 �yLT�u�C���$�}l�Fᩢr4����r�P�d
���t�����ڳ���pv������Ǝ�CL�_�o��׊,(wo�?�J���#��G'n�l�v��_��t��Zk�JE%��#�P�Y��2�-��A�AN/���|Y�Y����12�F~1��ӫ]��ӫG�*�^��7�J=�ӵ$\��#�':֏P��܀n�p�\ZZ241��L��O�,��L ��C\�]���SVnni��/{�d	�^�[�a/.���2Ԗb+�Gd妎���5�؉r�"Xq�0���a�rs��WI}>�Щ�0�6c�;s}�!V	�@����Y`"�vV�ۓe�\�����~R��������/(��`�}̨���>��7�L������ĉ&����.-��Bd��w��n`����+	\��`���+���A�����VSs��Is��� <�spP������ƒl/��l�z�j�uFd�;dn��ɸL��&��g/��ɶ8i���<1�ٚ~X�P{Qb�KD{�m0IU���S�R�~�UU�D"�pW�ã�J%_''{}|dXYY_ .^�����Z���4��\�s)̐A��,a�d%o�n���Ӂ�kTP��
e!L����M1
+�_ëZ�H���z��j�|H���t����a�wَ鈣Z���4F?O�Y2`�'ة�2|��7m�#j����M��g �Ŷp�ט���!�b��/���\^��,*t��	\*b@���鈝H��=+n����s;1��<;;"5�,�*h�lV5���=���LLǿo(0(�_{B�555��r<d�<����Y�6���I��Y���4bn��-c'�ȳSr�[�U���l�&,�a�1�vz�E���=��KIIĘ4�:�s��PS{`��Vh�^�M/PT�i���4���!4("�c���9�K�ƖjRjJ�0�����S�MX��f��?Z�](�j��*���z�sI0VC�yBȐB��'���������V/���zP=��;�堯�V�:g��7[�v8� ��^���V�ě~(h8ԠD'�ʵͬ_/i�ٗ�#,��k*}pT�����W�^�H���;e�G@���3!��[׭�*Ѣ���zzz �o'���Q�Us_
����kC"�� fZc�0��Oh��&o/�[c>���V��o���qݝ�ie�\@%�ɪ��}��9W�.����w��)I$��x��1�I�+u��\�����n�� �-A��{ˇ�?�0a�f,�uR0ǃ���Ta���-I&x�������[�ܟY�X
� E=L ���*���}�.�]� ���R/����~�٦ �Xa\a������$�n"<��їf�(3V"Vz���GC�{��rMlE��+Pi{�G#����f�uia��rԩ������^㕌�}W�[�d������'n�qs�$x�v��hf
�z�<-@�/w\
�1v9��=h�eg�=�F��,#8��J��4�x��v��k����P?�i0�2����ና]�D���Y�"�/�C�H)g��j���+=9���x���,<��4����,�� ;oU��t�`���m���`��ziZS�= �?��U�s�A�=��������L~�O�n@�(���l����cd�\���5U�˂�d���S֏�/�L����.�@���K�o���L�#�5�/���4�p�t�3ܦEk�8V�g����VC���|`���y�J2�*YS��&R�Ԟ�D�S�`u3���"��Z��m0�W=��mbc�z�X`�&��shel2��ļß����s2�5}�36�1����.��e|����ϳ��x,�Nn�f[��f��u6a���յ��R����`��88@�� pK�݅+ ���;��4��Vp����'`�Q����$փ%a��:D�$/��.)�d���nEn0�[%<o�.ic�\Ztˢ�z�p�(���h&E==���'y����a�A�Vrɬ�c���I�t� j	ʄa�XN.n��ڻ�ᩃ�0k���tUet5��0s
�m��b��MG�[N"�As�ڳ.*�6���NDl�w:_�w�y�]p̄i�7��P׃�f�Z�ؒ��f�إ��]Oӕ����G�����f,���+��&��sEH���ZEmc��R-3���X�^n?����OZ��Hl��?�8����e���m�L����e,Y�������eX]��i�n�n�p�71�C�}8�>�|��N˯���\iL�i ��4�䟼��G�U%�t�"x�6��{st�G]'��'�������u�1�`��@�p-��U99�SxD��{I(=������S$���`^��	�W_�1ǀ��F��-���f&��$T������}��Y�TJ����m�9�T'Z��9B�0}8�����e�����-�����W�S�yHqT/O؎h,u�i���h<���1֣�rM-�M��x'�g䰮7Z��:7�#�\s1���vE�W�����ǈ��	��	��;g���p%Fg�dD��X�u�� <�����1¾���M��!ĕML)a�� ��� āh�H}h�@d�ȋ�s���o�]>=;̜퓵�$���P�aB�늌qs]�mx8Ǵ�Ͼ^�<�g�P��,��7}���x�CK��_������)�6����~��$t�MB�3}�m������;~�	��|\��Y��ȏ�9vO�p���+d����ui�;�`�mґ�tDu����[$#l>c��^ʫ%��t'������8w��i[�t�HT^N����\�28J�����\=?|��fM
���>�Im ?�'�g��ȧ���z_��֓���(�Ubw_�U�5�^n���ʡL+�N�]i",E��NrVP�������k~V�`�D'����l��=w��gݜM��.��vy�X݉��(-+r��>���l���->���g��W�:?�i��a�k!0�}��Ʉڙscd�v���o����&�H�0F,�ٗ,�ǁ�����K;�40cZi��}0C�550���2MT�5�L���������o��C����Z�Y2�h����~�ۿ����ټ��9n*�5'�@���׼W�d�? PK   o�X<5P�F HL /   images/725e652d-7206-4b68-8c1c-12a8993f9b75.png��e[M�
<���������� �a������,�k�n�\���������c���U�ZU�*BIAQZJL�� ��WA���/HKaya0��X�Wc���NRڮ``H�>_FK���>>�ń� ��]�qߖ|��U���γ�Ώ��p��I�s=I(�-0;��7�:Z���%N��6�[F�w��25�6�eW��\0�gÿY	�A�N�"?L�)',�t�h��/,��kw���~+����Jad5�~��u��F
	K�"����������9�5,�������
���B��������B�_����V��؀_�����5����?40��ށ��\ʾbp�cL���9ߨq� @�_}����gS�vs�3s2����^l{\����TFLڠ��C�3�_|WD���6 �li�-�,�PXh_��`��Sa�г��O��u{h#�kS�.��$�Jh��)�f:�L������R����?|�ߘ�}��zj���5=t��ai�Z[�j�p9K)�xC�{��A��7�i��E���AQ�o�K����Z|쩣��J�M�Ԣ�=XJЏ���s#rl�����-�H>��6�\w��ZX홷�NyL�ӌ; ��@&��;��?��9��?������U���xx����[i���>d��f9�O<)�{��|nʩ�5ˠ�O\����Q���$�;i_n��_��qO�`/e���C��a�5�h�gb�B��	��Sf�$�g�����C��B7׭v��ʚ���0�#��Q���3��g�������!fc/F�[����r���^�4c��RM����:%M]����YY���ʻ<6�w6�d�'(j4��0�o�NX�C3���t�{w�5�q��j��%�N����z>X���T��g�D��<��l���ݟ*06��>��n.weeԗ8f4��0|i1_O����X+�w�9�����i�}���pWm�O��m�i}�GH�"�[��y�km�9y#�Z��}�3"�.ٗpm)�AעR<u��� 8J���Jr�K�w��0�߬ڔ��P�}+��P.4ְ{��I�����k|m|��/�����ǈ���-ϼ�'��U9D��&���ƬZ���6rg|\f5����Π�P�^.ܔ�|ײ��_�&u7���mѯ��-V׆�e9��VFJ�_�n<�OU��:*���]�����e�$E��W���+�xkeȴ.q�a���T<�7�P������X`Mc���g�{�mi{��f��:���Au�;�g��J�=B��}޲�I�� �3q�RĚ�<!��Pn��`����o�הGO8=D��M6ONHf��!�+1�"��K�������h�u��S�����zN�QkW��~�זyv�-�4aO�=�8�f�}��P�e��4�X����C������.��h�5�ʃ�����0� �)�)&oޗu-p҃��zl���g�+ۇ�>��0�̃D=�����'�>����5V�G+{&��+����������+��ަ�:�S�a�45s��ވ�.mfK^j����Ǌ�f�5��Z�)ט�j������RM�.�BȉLq��S���wߓ���R'�q�cuZ�s�&;�[ @�X�o���]�W�=SmI(o�e��]$����g'zŶh�z��>Ġ)����
���R�o�h���><"a��f����.��{RE�2k2�d�Yg!Epj�/���hC?O����	z~�w�����}����`�~Z�L��~��,G��4e��?}��{/��hs�����i^�դ�P:�*hR,�JD��]d��2"B���Ͽvz�Fwz�H�$K��#��kgc=��d�n:j?���u9�J�v(�~E!1����;n;K�zD�z"���Ɩ�F�{�Lw j��V@8-�B�|K�4�A9���i/��m��1�� ��xju��.L�t�Z��Q4���H���L��m��P���a�D�T�DO~�S�~(Z��IR��;m�N4�/q�.�r@��j��3�F8���?�Yjw4l9�鯝�M	 ��}�?�\��f�*�U�8]���w?��Ⴒ����x�%�ps��U��i�Aɜ�x��s
�!�$D�^9P�v#yE����n������K]�&T�7�at��]i"�R�R�ҟ����1Fz�O�GJ�n��9����C?*w'>|��K��/�@44�#+М�AA}��BƾDZ���b	ńJ l���l���X>1�� D f���Q�aڌː)m� a��|���%�jJ(B2�v)ID�Up�,{	��B�_��ܳ�o�?�@���<�M������\aV��oM�	���@dx�c��0��4uV���N�B� �y���� ���q��7� UZ�Z��L��^Z��{�(Q*�wH����^�D.O��S(�N�K<6i��1�B�"��<:z<�u�J�X�i~��5"���8�e�}���L��f���7&� f��^a'��nr�5�ȑ���x��#Z�F6]fwV��{�O��V�b[�<�jz�hE�0b�E�� �ݼ5��WH����}�]vͬRD���)=viĦ���fp�#s��OO��<�j
y#��o��c�`�K���*.9��{��Ƃ����9J}�cx�<(͝�{Q+ۛ�L�/uuT$���dT�?=�"�{Ք]�~��4N��y������ºAS���onܮ �?����"U���5����!��@��ⰅUrO!
�A�"�����)��
���h)��tQ���KBՖ��[������1�ԇ�%�M����W�m�4���{���O�ȈLwئ� �_���n��vօH4$��-+/���!͟<��"�à;�����uj�+LuF	9���t�u��D�Ų���꾕��~�,9��Z@�V�߉�RA(��"���݉�V�S��F��t�g��N��}JW�G=/S�����Y�q�熳\>d[p������I*]� Q��,��mF��>E$�\���)e��G��_�G�2g�]���T�5��$���V�Q�
�o�R�;w�ӺD�*���v����>��$
Hu�O�Mr\�c���Z|�g ��~������w�}h�k��*Y+�����pНΓP�'i�����stq��O���*��$��$�j@�Z2~�A��&����vM8��������a�K��/�I��!Ɋt��C�EV��WG�L��Qv"������iՌG�ᣔ�-��=�;�90��� �Tv���^�O����s���9�d���/ˤ֭���!5U�S%��g����ťC� {P�ۤ�I�)�3��G��?_������|����U
�}ynR�s)P�Н���8$1���¦�2W�������Q İ�'�؄�F��.@掴��F?<,�L2�8vX�f�������&jk�}����I��ʒ{���T7o0Z<l��XX7Kb���,/B�g���
�ʿ�)ïz]�{|q��3�T�����=ӸUR7��4s�O�̰�{�n��t�j�Ur�I������|����S�G�w��t���"�g�o�7���'vXC�K�Y5����::km)㥖Z��hL�ӍF��7� ��|d���`�8�s�j����{��IՆ�W^>�b��ib�tU�'˭n�Ҏn��'��_S�m��J~�O�|'�.IU�jS��׃�ڤ�b0�
P����^&��a4�߆ț&s>#�sc�a	�[�]P�I��0"'�����x*�Ӹ})���Y����c��/�x�/����*�Y�̼��Tt�l���jg�/I6�Q�i���J��Hp]#nߤ�&%�ո�m]W���-���e�ׄ:0ZI���ˏ.��%��96D�a��i������@���)�׳G,��ߪ>~���-�r�*�U���{����
q��D����{��~��X����ĉ�p��s��_�t��I~�$�eN�/P�Z�7Ue糱��ٽ�g�U�����^��J�V�)J��B�<~d��[3ϑAd�d��F����$π�'�Gèpn,9o$jd[d����І^��}S�T�͉���x������i}�aFޫ�槙��3��Zn��(����8���C"���!��.�h��� ޼0J��˝ߢ c7��8�/7Y�)A��%b8��)W�o\,�4o/_��kJ����`sx7B��I2',�\)�7;�r����,�Y��-x��p��Q�`���^,���jb�,���PWef�+�y�`����c��i}>n�g�u��zP�pM􌓐a�3����*U�d���[��Za�%�ע �}fӟh�f��)���tO4s�:�߰1�a0�r��'<��D�!�+K8H�t'��;����Ѣ��͗���x��\���%���:�����1���̐-͵��!G֓�=�!P8��*t�0��D=��<��A:����R�ݷ�L�N����D�:�N��_�ɛR���=�=�·�
��b��ڣ�IG�~T���o����l����m�����i�"I���H�*���D[�B�\��D��&D&���i��D
��U*U���U�����k�K8n��\��M�mV,�{Cо��8�����H�u�l�صF��6��MG���-���U�68衂�SU.:T�j�K�L�ʂ��93��L�J ������ڛ�s�ڋ�� v�M�D-�:���y���Γ��h�f{�fb����.������u�2�i�����T�TM�"~W�O�x�AY��v���*\��
� %�՘��O�6���j֧�-�ؑX���=�	:�&	������XD��a��\�m��~�)�p~3�(8u�`���X��dr��x��y(͜���ck-�7Y���S����Zzw ������W�Z���Ѭ��k�c��>N���Tf@K�T4��qv*����\�tX
���( ��OǺ��'G��a�x.q8�:NC��`K4�4,D:h�L���`F��.{rk�j��9��4L�� G���Q�(��{>_�/���a&�v���:�e���8��jZ_�O�W-�����N��Bf�(S��/tiT~ޡ��2ْY����y����1+ѳ�s��d6I��+��o����v��˂E�K;�#,�"6~8}��y�wb��edd�8�����?$���cv�\,���h����L��zj�����&�Z̔�%��1Q���Ns�i9ȏU]�Ō���")�+˘�9v�9��eeѝߌ��)#��K���1E�	�`yu/jȄ���t\���&I�B�y�(Q�XoB�C`��7�|��rT&_��������eLRX�ۧz@Q��������뒧+�3�l$a���
,��n���b�m���t�x�0Y^n����o�_��<��}��Ixk]�����;=X!OO�Ygy�=�qp?���3��H���{3�b��uw�`V��Yk-� ���($<���4�4���Z͜�1����5>���ƺ�M�UC�9��`FG�l�|�m&#ě����O=�A�;O4���q}�Z��0��#M�F�U���]u�ɪÊ��O�8�͋.O�&}�9�r�;��1$��i�Rq]�y��Tݨ���F�6�Udtt����+2���X*.3������� kC��X�;n��m���{��.9M"�l�g;������>+� ��������Bn���f�ΰ���bG�{��dc��~��k=LM ��$�^��6�C����fn���щ���p��kY�.6��$5��z#�@9s�"�)�!��̛��,E�}�hgj��ۗ*�ړ'��1 @�ʮ%T�dG��kٲ��ֲݹ���tD�����vQ��F��6,�����ϐf��I�Xn^:����3Aw���5��7K���=��_5{��Z����q�7�um�:a����2�/2)Mc�8���?����i�^��ME�P9�_'�������B�Q�{{_�9��{V�t�~jI� �{��_�ZBxz;�}CY���S� �'S<C_G(NW���d�+Q���a�։��<����#��yJ2ÏS?��K�{��Fj�6jx�r��;�j|��Bҏɼ"�Xb롶���&Zy\=l��切=��qL��(�n}��Z���i�ǹ�bl��5�N��]��c���AZ�V������H$��|��(��}���4*�(a���Z-l�	S�	yَ����sl��lh�fg��^��4��ഏw[]�ݡ�q�-K���Bgafv% {D'	I[�?uu�՘~*���U��٪�t�D�d*�~��� ��[��;�;a�n��`}6�4E������_��O�>Uɻu��H�ϑ|I�rTR,>i�P��߸���� �x#��*�I9�:��E��T�'����)��å���Hnh�b/�����Q�l����^����q	�+.�������Q�V1ۿ�[a��VR(��
^�L���x"1x��[P��-@��#��3Ϋ;I�62}d�&Q�i^��`����;&Z]3��~�%�A��{2	㐢0w�Pܰ�7�aĖ��2Jm���>�娵iQ��E��ߨ�l�b���0)��o��%�k��RW ��/6W��M�
��8��d�����/3�2�wY����N�W׃�qV6�Y,��0Dr��5��S� �-�#t�����rI���{ǐ��� \k��	�T�J:A�B�0���A���� ��� �Ł�_t�G:dQ;��L����=�����t�x�����_�D`��.�ďcx<��t�_	�f���&s���I��1�x�@;��Q1�2���D���Ŋ�f1�A�G��F�jC�$�b��3 ���_�1u�`��@�[�kJ~�\Y�A��_�h$U�`v���Ip�]qo�F�f�/P4U�¬1����:�Q�#t.85u�S����v�k��Tlq��L��p���n�(<��z�����ZUkz<sJB\��I�؝.���?�6cu�G���0�,�ֲ��Ɲ�]1�8�R��Fg�އ")�Ӈ+Xu[���a�Tf���\۝�V� ���F������$T���Q��w����U�oK x��Ӌ�����x�E�s;�8�B\�4�E�[��Do�Qc��6�	��ۿ(�`9`��{4��/�>�\��N���E�uM�Clz��8������7o\����ۑ
�s���k:"> ������,F�N8��$:7��=�r(��Ċq,�w������v��YO$�1-{J69�������1�;k�'��-��V�B��s]S1·'i�1^��!��"�R�,R�iN���jhp� ��s�M�p��1>�̳���~��y*ң�<N�����������n�������kd�sqmu�`�c��h-�M/!�YL���ah�p:;Va�6��j+�:��ƞ� ��*��T�A����q{�r�s�a��P�/��}��}�xnQ��o�I(��Z~lLsv�qHG���I�Ո����;=�'�ٚA�Y]Sf�ɕ��L�3����Ȁ�T��Tp7.�W���=*�EV��?N��?n�W;� #��@[g;]��ҷ�������Ă�i�\���#�~��{������ʽcXb�cњLy���A!"��ݤ��Ts�S�)nǣ^I'��]�����p	&w ^��9&k��+�,i�7�DѠ¨�T@{ KkՍH̯�e��VT���"2�����i�}�iGz����S��ߗ2��\�#r����v�}h�x�;v�!A�@O0�Ar��p��0�5D��0�����ү%@�⁰�d���
|Dn@��WU{��.
eɟKF��֯�����Y��7�=�ӄ���H�"��'����3S{ǝ�6��i��u���y�|.�c�T�����)ئa�\���j��k��'������ֹ���(Qh�TQ�T A�+�����w�mS��� ߪ���病��s�2a���t�����D*�2-XnL�ߤ�&��3Ś�h^~�Փ��u!b�.�@	� ��Jޑ��QoZB�c�d�eH��O��F	������N�3>g�X/5�YUUj@��c�W�k[v8l�/��$�������P�d�e�%�H�����л<��{3���|��B��^F�pa*��A�w�Q%V�!���\C�<�Y��(�{X�_r#X����e �m��qͲ����UʵfB*�P�d(�oE�䠱4���������WUɫ!Io�� �X�?4�d����f$��<�ǭ��GE��~C��Z�Ș�#:�v����:,H6�Sl2���.u��I_};,����$&��H"/6!n�F����5!�3�Q�irDtm@�q���$Οd�ԟ���z�d���S+^T��M.]e�C�Bi�|2�)��_Q��oZ��+Nq�lWZ�D)��r��x!$��(p�N�h���5=�T
�}�oV�S q�Hӕ�· ?���GA����D�����t�w�ߣ�����t���f��!������a�X%!��;-O����:fo�@�j:9����%�`k�`G[��'�ʂ��ɢ^/�$3�_��e���<[*��]DP(�VR��w�\}�<���{�B�@��l|�$aV��_Y�S��!��D��:-�����P���x�31�����c?_BǍ˝���GG7X�ۗ���%R���KC����܃h���fƩ�{���g��6�N,��r�-?^:�u����&>���?�Ff��)<X��]�}�7�I�����Mx�hHЧ�?e�9�2V}↾�/P[����TjY�������p�ya._6W]F�R�����Td�ˋ��T�%99�g�WbD���8�z�����"h�����q�
2�@!V���Z�.�-D�ۜ�D� �g���BP�a�+��e"s7� �Mx~AM&1�}���`Z��@���N�����ŜQ��]��<24��rU�����&2bI��]�55����Β<d�6����8�.������	P��˥���.��l����4�{f�2�<f�7T�=@u��N�a3�>JU؊�CK�M��I+9䩌�������	>��*L�A�%1Ȋ-�*��u�qC��&���i�������sgLX� ��T�S�Rc��HX��2�t~= /��D���
J�[}Y�
P��#l���iH�*ULyS�0HP�4��:BQ���'A����C��C�K����ҫ�wO�wN��,���fRu�L&9�Ao�W��sf������]��Lk�g%���Y���S{����Tk]\[�}i�j�F�aej��R�B��W�W#�b��s��P����Y�(�g p����,��ur���%�y��6�*�x��O�����0$؏�S��u��0�� ��嚿4�ށ�1"e�u����h9?��`|d��Ms��.F�J12N0	��q�U��,�#	�5O�� �c�^rzP�Vh���U�mz�!-aծH��҅��u�@�fH�ݤ.�S:cc{y��.��k3�Gn�d�|L�k�߇D:&��l�����G�8�WM��<֬_�������<�}_���#�^�*�0念4?N%��K��}��<���Ē��E0[`�Fh�w�k�ٵ#><@i�eW�p�q������~���Y���?uYw5����G_���e�d�c�b�=��Nt[�~��5��>��_�MÒ�Z�	�|���鍦����}I �ќT|b9��"B~�w��ٌƇ��?[)�YQ�'��Z5�@1'8�T�.�]��@x�#��*pFwn�p�$:�ܛ�sp���������<Ww�Y�'���/-���#O��qf���6G��+x����F��|!��5ӱ�C�D̚�D�d�/>7IY�s��M��<,�@^�sX��q��[�H<���xE�����u�n-�̑��6��tbEB����N��N�u�S{�L�G�.�L�""Мj�F��`$H��.�̚�������A�A�}��s�<�v��&S��<�J���(]XL�F%�6`	��<_#ȼų6#Mr�&5�@�c���E������R5���W[YY��`�ௌ�4��*/#��Kh��J�ބ�竴=�J���N'F�+z��+���!��]+|hp�L��WGwBA��mH��*����Ny�Nj�Z��{���V���˃wѢ8�?nH����M
�SV5���;�
�Z~�/s�٠�w�f�zq@��_�Qn�Hn��{��6��m� �/��J=!z�o<�u?T�C���o^��q+F�)�'���^ ќ�u�:�$>UL��B �Ճ�]��ӿ?K��C<)�c�F���V7�;;P��f�D�+�i%�v
JB/�"� �[�S�������N~�a8����*�I#���&栉��N��-�l~���NU���NXB����'v6�񀧣Ώ���A�1x����EB��ˏ���]�Qx:V�����c�TK��K��ѹa������)6�mj�o�I�ȸBY�'�J^12�KMK�=�yD�ZLI9�(䣭n�e���
�B�
#� ���^������B�^����\%ᜇ��9�I�]	4���(l~��YI �y��%=�7��3�h e�q���6��v�����Y��@_'Dh�tW�����3oDWk�S�����cD[�R�O(�,�q�:�J�/͛i�I_�&�c��98��(�\;ji?���E�B�G0��ĵ��,�/��9 n[���誸����Wt�פ�E�׋-J���.~~+sU� �=�RD��V�S`���#>8n6qn������P�>�C$�pA���'`Ga���l�%�ݔ���2Uqq�G������r�Y���U�le�1L�=y�q6� ��-�S�����](xPejďџ��[������q�'�5�.e����7"	1����Q`Ah�u����wO-!	��č�k����L)�q�?����\�/�"z��u�Mc(/�'��d��|��J���<T�4ixqqaȊ0��^<m����$�}絓�2_ub͔�Z;�lR��(,�c5��XYɵ����3�P�
����;_I[}������+u�ȅ߈��Ff�a4�j�σ�q�R3�XT�d
��N|QS����ꌎ��O���Wހ��j䦄w��7����� �I��{'��w;GQp5P#-L�"�n�u���VvRy]��
�3ﾊU�w'�8�*�&��ԑ�Sq�gD�j����(f��t�І��嗉�*Ҥ��ߎ^(c�\U�~�O�ݥ�=M��E���<@v���A���E~P�E�F�e7
J��K̅�7`o����w����LD�0�X���d]�I!�$��U����<��*�	��T~g�����Շ���"P{�_S�>t����!���2f��phb����%�TZ^�
��*�l r߾�p
7����
<��~7���X��[5ضloO
9�n�F�reE��;Į��^=p�0pr#�  x��Mt;b�,(lgog�k��UU5���5!!\� ��Vmf4�����T9�0�S��:To�.Ĝ� ��ĽF@:���ٕ?��y|Q�6_S�8D��j�M(����^l�B�uYaU�X���/�mS�镵U�Y9�)�:a���5��P�;�qr������ ��]��.�Y(�c�;���"4����nOX ��:3�0�P��Y�i�a�b�V�����[������`�4ӮښO��4�4�9��3@��$�(�~S��O� �^�a``��`f� �X�b��dm�ǞtM�`���%A����!?�{|�K�Y�����ڮ��NN�y���x�iZ���%o+�/b�=9j��2�?�EƮn�5G�.����]��Vɑ�.��x���`,j4.GN_��[3ɣ�:-fc,�����E��]3�R�n�������s�Z�z}��-|��g���8
��[��FIa~/z`Ld��eh�'�ٯG~�qGf��J3��ap�$ʫ��rtض��n֯@w�K5��zl�Z�'WY�H+�ZGa�NGkd���슙��v��,�|#\H"�:�-`��aל+^.��ꂏ��������fa�=���l� ӡl��p�u�q��m,D�FeM�m͉ю�8�
�.�F�7��,=A�� bArj�9�%3�m�J���M��cyc�Ki�_�yi�p8�5>&�������>�\7��G�:>L�S%�\'�s��&�;+�G��4#x Ir�gq`��@��d���T�^[�'t�&ӧ�7��J���kZ��:���PZ_u4�>����P��.>L��u�V�����:��H��>Nٝ/�UQCK��q�����p�;V�����6s�^�h�7sUK�)�U6M\a�~.�OB��%/���f`�Pcˬ�^��
�=s��l�I��I�#%1}� ��	`�&T#�E���ΧLR��Ӳf��C3�\�Q�z�a�Z"�F���/�t^&s����2�?K����Q�^Ө�]��\(#d^2sj:u���z�	
�m����N2#��G�{֋��������������?*g��J��ǜG#�����)���[>Uvh{��=Vt��j*�ˬ=R�WU���8��6z]����V�h^v���cUF7¶hZ2�}�l���0�x�6��Hд9ձ��ap�Gi��t�4�u�E�k�!��X*�!ڛ"�XڰK�IM$%��N?;B�(��D-�X��O0F6ە���(8��V�A�n�tӗpJ�\OQp�R��2MM��P�<<
*W�Ӹ��Z?as�g�� zk���|�m| ���e�!{�Љ�i���hF�ٍ�܃xU��ⵯ�ҽ8�ݚ:���y��&"r&e\��YW��K���8�D2��l;'��/Nf�;=�:�i��� �OBl�����S�y�~��i*o�$7�Ἵ����Q�ƣ�+�r�b�x-n��?��Û����E�<����m*\.w����'�06����<si�o̥jUJ���\���z�~��p'��P�����]�Wͪ�d����S�}0���(�-��-~�'c�4�g�@�
�V���Ǟ������F%�w�u�0d~q1j��qN��_�ke��Y!�=iC��I�X�B���IsЕn×�/~���Flb���"��y�9�Qr��&�J�=8��Ð�-�<JA�+����l����������ҤR�h�ϲ%E��{�H���T�����q��]i��H%�؏���,2It2n�dvq�]u��lTZ���n������C�'�����!ER�{�8f}z^Pp�wQ�{~����y�5�Ho:��%,0�m���h�8P��������S[����91w�g�d[Sh�fv�O�Pڑ<���_	�-�N���k�������@t��܁'���#��~��Sh;}&��n'�E�|�D�T�*']�;ZZ3� q��qn5�4Uۀ�<���C��c�ڔ�#'jL�����E���%������%���P�
mw]� ��wwʵ�0�D�)105l�M
bɽ�MÉy�Fp�iH��$���*ĥ�_�귌�f�+4�D�|��� �E�=���4�������1���v�Ǌ���h$V�]� K� �'憩(��>'����޹K��'V�-�2�'����������P-A��!�����)��89����Y�|���ri��av�D�̫�����RЌ�q�o� &ӡb4�}��v�ԋ��&�Z�D�)�~�
8�.��}	Bz�ȝ8�����Yb����u) ��z�ҲZ�%�̏oUG%~{f�����GQ)�tܥ�go�����Y����詖����4p�a���C���I�������0Wax�J�Y�ϡ��!Ґ�E�X���`�e�;]7<�0?P'h=�����p�.c�rۦ��878W*A����_Zz���5��.�"KP<揨��m]H������',�WD�t�P\��y�`	�5�I�fb�� ��ڋ�)fw�uF�k�KmW�<e�!(@`$x8�Ǐ]?���޲K��$R��)�EݜUYFi��@;����z�������Κ�����ɮ�����#lY������.�Y}�_	�l��h;�@q���~�%��>HV�.�3��2[j��mq,j��",e�����: Cv�h1�U�E{��ņ8g6Xn���Tyy�5XfV"��elQ�h��}��_bQ6�b_��f�Ms���o)���.��n�C�@3y/��F���0���� sb��r�ǀ,x�����7*�cb�75��(&���������`�_̟�GY6��9������Nx+b:�����s
t�`�\��L�Ӭ��(��q:�q'�������._BZ�����ѱ����U���Œ�V��C�X��"^���̆����G=��>DᥥN�͸�<,it���?���_������^��a:�WB�=n���g.w��.{�N�:�WjI�Ku�q�Eݭ�%�/"i\���[����<t��f�YȗH�A�߲�F�x�K����V3�U0���L�%�(p�Ѭg�G�P�,%��J�S��#�4g+|x�^��[w ֹІ^������j�"/)fq݌��?t^X�������M�62�?1~b����81� �vz|-#������io�ȇ����XX�i�!:��t}�xk��j�vw-3r&_⠙%_��[Q*|�4�g��y�ɷ@0݆��i��{.NT po��p놯�̋���o*��Ύ��&���(M�6%��#8>��/�UZ��,Ť$��hQ������ț!�3��ђJ
�x/o�C�|ݡ��������|�"b�+���K��Q8�W
e$�����Y4�hE����+�.˴x�A~e8X��DS	G���L&D��#-4�IRÜĊ��vZ�Šp$W8��z���a-ŇW��`Ɂ�i+I�5ӝ���u�k�B�AM���� D�i4թ�����4���4ls��9�P�^*�<O�Y�"�G�2�J	S�Wl��\*Hꂱ�D�v9�p�8q��u0Н��?���Sv��!�O@.�o�U����1���!@Ǿ���E�]��$L����^�VA�4�kD���4T�3<��d�l4�8�4��0��umM{ʫ�.�^�(B�]ػ���M�� �;�-M9�;jZW �
�C�Ē^?b��+�,Bp��@ @^�ć�����s8�����2����_2��у�9˾�@*Aa;�H�M�k�X������<P�ǴL�,5�8����#e������gd�Zpи����Hu�q�>�j����BI2��T�>\{�l��Xp��Q�l,'@AS�C�%]0=88w������j��]���������_7�<I�M�;w��?��r�"��;�#=����|��v�,;w}��^��}8���g�۔ZV{ql�Tz�`���e$Z�E�}V^հ�dx���|p�F��W����/����Hӯ��5(�c��}�g��p�Z���FLr��
X�.�����q��O���e%G<�L�)C1-3����\�Ƽ��jG!KM�۹3�t�ʉmޓj/yp\�_��C�dN)�<�OYIA4�a�;��������Bh����T�']��]c�:��,^~��fN���\��|;�Lr#��)[��Vy���Q�hgyS�,��֔c�j�v;�ݹ��<�#�۸%��?�����z �}���Mk�]�͸���pVV.f#c�)�8�G�7x�L��3�
��2��ѯs�(�6��*����k@K��P��Kۘ�fzl��NZ��q����4z�¾�`y�$X��)�V��v�j]	qQ�����E�wV�R���e�ES�$kz��H��1��ކ��D�w�+��7D�DE���{��b�.���w�$ �Q���k0����E���>�6J;dYO�k
�T{�m
7��%��C55���"8�	]�ј�񖽘��w!;�}��e$���D$����!����t�D�.\p�qW�wVr{�#�#��!����}φWQd���E������~�fC�s����6���߈1\�3fص�c�����'F�����V$G�kx����v���o�d��m��m��I��f��A=�����͍�D��� �^�A���w��`�m�?9� Ҳ��|("���[���M/� ����q��Lڀ���Ph�8���4,W�""�+?�)�AX-�#�݊�?O".zBFCbג�h�W���_̐�rj��nL�ɣFm`/�v��;0�D��c|������v��y�l�j \Q��#�����ѭ?�.�r����2*��i;	��������$��,�%XpwwBpwww�������s�LOu�%��}�� �z�6��tR�|�&���	`�ȃ���l<�'{?*M���Id����nح�6�!��Y�r��ʌa��b������!-�X ��l�Lx��u+��퀺j�߱�bnhl}]ZZ)�����p��K�
'i�3���d��uץ߈�bLI�BU������nW)�&I����5�B�{N�����5E��#=��}Q�#��u�u�O{�O]#��ܯߦ�����ǽo��-�� �ǒ��]'���I�w.
�jG�ֺ��`)�cH4�Nf�mbb,ZfBcbDފ��\9_�=f �[��g���%ZU�����$n_Fa��g�P�6|�1o~9]`k#�q����5�M;��h��?�H���9�*3<N������6�J��s
�������'Q ���m�闗������ת���PLn��
WK8�`�G��>�%IƯD��)�r���*�\�1��;O�aT��OBx��i�V���n�
��΄��F�Yr|� �Z�?�J���9#y�(�@�o������$u�������?�m��t# ���!,P@�2�3�nch�c����A���m{8�Y��� ~`Gn�a�K8����Bu#��b��@�͙9Ro���S��{��3�*X�m����]�ӉF�rbaݢ��������Kf
X�k��;�b��z�Z*�6��A��7>B#��8"o���G�1���YM��I���3�4������\�9�"����F�b�����9��{<�����t�iI��S/�����p��n\��>��!��p<��e�������Ƀ���wk~T.�k�Z�	��t�g��d���:�j|�X�\mFL�oQ��O�L�~���TS����X��i�石O�y{8� ���~76p��E�����ybn�ӯ��<~���<g�S���,�P<P�]+�@F�I}/jq[�B)>g��o�j�rs���P������Z74���;��Xn��&��Y��Ob��v�k���)�%Y<�݄���@��+���ri9�ɩ�1k>~9!e��ep�*0���R��7������NA���l#�*����l�i��vw���c���==b���i��.��j��k�e��J���O�z�Fi� ,�����###`��-������/��1M�	����]��U�Fen�}�~��[a�U�hl�r���tl�c{{�@A��o-V����������=N8��g����H���կ�u��6��T��/1++0H�����0�^3?[��H7���4����q��OV���Y�����+���ڔ���KG�&�^�R �����ͼp��$QYы6ٛ�Ӭ)`߂p���Xc�BM��,'�f��}������`�m�6e��h�#=�l���Y��[�6wOC����US����N_w�6�~ׁq����Ƙ���e���b�~_T�®D�W���9+=��h��'�t`j�^���0�9�[U��joW�#��u*��n����q-R�� �R"3�W�
���
*��3�񲂢>�S�:��I����Y(���?b4y�r糭���8��l\���ÛN������[n�mH З�9R�iwB 8������{o(&�~���|���yѽ��q$e,�ڴ�k�:�>/��*)������0��s˫�ů��'��s��M�YH]&p6R��t<��b�	5��]Ucwt%����^1�0��b��2����m���F�h�`�:��b~�45]�8#0��_��lx��Q�خ�	�H�J�HpR�yө�ξTW���S��������aڹFy�r}4T�b�YT�|4�G��_mKTWJۧK�H,���(싎S�}1����κR�RX5�G�\�k����c�*��,��Qywh���(V�&�]����Ǝӳ����LվS<��=�.����џn��!Wٱj�=�|D^�8��>�>u���~����um�q�䇔-�cbmE&���i��d���w�>&����=�@����k������������������/e&Vx�O%��($e��P����O�¢�y���4���3����3pGs�Qz����O@(�dI��u	������1<����y��SQ���y�')�xB<�j�!��O�=�A��(~,�`�����6ޛ|���X:.&�:� �u��}��B:}�:�+�}���a�������q��/I'���9A?��I߻���2��
�d31�n�����k�JDt��s�Y�&Qc���4�rjyU������).{'X"ES(G<�\c���Xd6Q7;�a_V�1�O�*\�>�<��)U��+���9���q�M���[�*:4ɔb�zR%��*ʖ�˰ˬB���r���(�s6�*Y~5&��I%G}���ĺ- $'�fo��n�㳇-�.��#��ݐ&k�?�i�_���kL	�`�Q���(�[1CuEc�4��p�6���Z�Il�݂C�@?����`����E`�	����2������~�c�Ei-�%�[�f������Gt��+����M&��m�gp��fx4��90��'��Z��d`O�d��s��o�ڨ�i���05�>6#�E�L�:�#J�fM{>%XX�uV|���J4�W��VT�\���$=��,���-�T�.�wd�Sn
.�:mX����S=�w\�FL�'�My��L��R�"���'��2�D��*�l�f�s��T"�\���[B1���$�4&������_K��n��CWݏ�w5���>�ֵ��ȷ�'Y��ӏ��5����&j��ż��˩��(�'�N�*G'��B�/�sb�Fm��ӷ�K�9B������{���-�ף�����owˮ�������D�1Dw>V�Nb�������%~m�8S$��Π`G�ҙ3YKR>�j�5���(2��ŉ5�e�Ȅ�"}�����tmК�_ bNe��:��2���	Ð�1;D�H�����ߍ�#jY�ne�x�ds�W����0gKI�#t�?��'h�j�����nҔM�N��䒰��_F��y�C�2dl֏�E��%���۔�����1R����#�6�M<Zn�b�8����m^�>挗��P����/RY/���b�!�z����uv-m��l���� ]@>��?��A6����E"��:i ���w�Cލ�)��ߟ l!KTX!�s��M��d1�$f6����0���ְ`KSxJ:�=�'����Dg:V�v�10�>8z�x~'Z�ا�WP�M�<Xt�fq)�dx��|3R)(1mƹ>��gV���>ȝ˃8��ט]��\A<��ճq��IH�>j�-,��[�@��̆E`��`-�d��s�m�,[���@A��B��Z��1�,y��ۃ{z�u}��q���8
N�t��,82�������.�pgR	F����M���w�s�m��&8�f��Q��f:;�����F�?���L$L;�~l]Tl8�Z�E	P�fZ��(�|ϐ��3	����P��c�ї�7!��v�E!���t�	N���&��r���ɼ'�P��u#5� ��ġ���kX# ���i��@�/q�"HH�*ߚ���n��u�f ��FV��q��$��i���NҀ��h�������h��/ڛ�D#��yª�UV�<{Y3PW�S���롊��۠�KaВB\�
�:i#��p߫�:N��b�l_�|%�V#&�f���	5j�#���V�%(R͸U�V�8�w��YG��5�1�B���+�ϴ�_*M7��=.���%�!�t���qj��T�J^���g���Wl�����Z��(�h�9��
�x��8���*��V�׵��i���W%� �X)���8ln�HMv
\:�𮸪'
���ϓѹ���̦���U��ސ�9�st�h��^Ku��FN�ǚ�L>;�����%�h��.*�c��h6�Xuw�e]�~6�9{PU�?�B���O�]���W�5�l�"EµE�(0+U�?��`�0Z�o���_�Q��G�\��,4u/osƇ�����v��U��=��fGS�JM��m|9��@�8GHO�ֺ����]ot��	���2#�l����$���l�w0;0`�Z�Uu�*���V�q��GZC��C�a�`�rN:hc��Vi����g�����_L��K��Z�E$xYݤ�?���@��\���J������V��ղ`9�o�Kd��H��~��N���cO�<HT��̺�-�b۩��{�O�J"� hX���51����/E(�����Q��֠�ď�`(J$�\���b�t�8M�c�W!��Oz/L�<)�]� ʺ|�]�ik3��1�o�����qA�`�ª8�w���q%�ʗC`�\,/���q��NC�Ñ
�n6D�U�ڰy���_C�w��f����$ Wy��To��<!�(���΋�(Ô����)�Z5�W�hK�%�yZ���54��Y�&/�p��?7�WGv�u@;�0�>�.$�����|V��]:�l7H��/�#Үv)�O�}(����~��ká"H�o���v��CO�Oc(��V�e
��Sm����Hg�j�(�L�{�ɿ,N0�Ǉ.���zQ*CC�w�D�fg2,�L�K��;��r{(&/�!rZ��1�K�AU� Sk�&.����f��>�glO�����j_������l1�.�Q�-��M��l33�b��6@sg:���q��(*�A��D��N��J&� N��Z�Z;�摤�@�#��ڡ<
����8ZN-�:��(0�W���e�"E����'0����#��Ol�N2�����:"��af��g馯	RX?�z��I����Ah��|s�F�z���q�ǿR�@��.�BڙJJ��m?��,o���rR�V�SPBH5��R<���z)����=
��Gcp�|�����,�zVz�+�Bh�7dj���/WE;���]W�2 �\N����2jS���_@˥��b�eOo�r�Aw��4-�l�;x��;$�&��`hى�J�)"H梕>crs'I��.D�M�zv�?�c� �"ä8����Q4ԯ���X�~#T~؎u��0��tg�P�v�VG�=�Էم˭�h(���W���e�C[^��|���٬� PW�f�zÐn8%T��O\���T�|�!�r��/��"�~�s���+��OK��������b���n�E���A�ˌ�dw��̍�'�۾�s��ih5'�1�I��lLyAI����ᖶ���1�&ty���Ra�d���:��~5ofHޣ�y"r�Ta�a,~V1MB]D����8���ꔿ�X{���g")Q	8� Y p�		4B�O�P��MQ�/˙���!RIΑf��/-�.�B��2��m~r)�/��׬�|\G��.����1i��AB
��ӳx��e�~�.G�}�ʲ|�#��$>��l��7U�N��E�ٵA���G�.*Rv����zW��,@��y|����l���~k���l�>��"���T�&un�|j��w�{�ȁ�3"+\3��"r��ރ�jIh��H��1d��?����j���V0�%�gZ���;����5�n�� E���-W���=��U̗͛��	��K4�g�ǵ�J�Ly�}r0�89��� ��e)�3hhYb�%O��Xf�i�����o��$�h��^'7>SS�RA*�DΕ�(�3�=������'����hbm�������TPE���C�3��U��\�h{p`%cHm�ecJ�u��F��R����kH�e>VX�I�{�c�M4���'ʆ�4�#�'���|����!Z� �bs�;��~�l1�p>!�j�B�f������I�D��I�cE!�F�g�ޮʟ~��M��$Ґ��0ݚc��$��3��%�t��5f��b����>���k:#�&(�}8�qp0&-%m�}r*EUY���ʕ������A𲗇�������p� �[	��&��_�a�6�-��ڹ�m5���m��ޘq�F���@��W�6!����8����-�����l�	Ĺ5��ka�W���*eTď���l�y�@��V��H�{7���f�R�8B̠0��s\t���z�Ŏ���w����ޮ�?9Bls0+��\f�̈́���s4�\�Tl�6��m@2�����d����[�QXw��_0~��^�?��������U�UC�3b�8Q�q}.]x#�u��&�����V��C1\�w�I!�	�RuT5����㶟!��ll~�@�j�zhNe_��(L( ��V�� c�;��
'B�iI�w�D��-��{�X^��κV�`6�!��=�g�>���-��]��ӕ}RNR�wm�|al���W���KR8g��P���/�z�-�¼�:_��z5\I�pd��M���40��R0˶��rB\+[��fh���mD�9�����җ���W�$����=Xi9�9�G}���E�6�B��;\��(F�]�G��N�G���+��6rD�\C��~��al��T�2����P;��)�7�9����/U�ذc�d{�����_0�j?�ؾ�<u�%��"�����=3����U(�6��#���o-�R�4v��h�ģ՛F|�dEJ/�hBɲ�J5��pܼ�B�o�sp�K�{��_d�j	��=�Z&���p��6C��O�c���Vz��t�������Ң����s����)�f'Ae202P�/׽O);��������M�s��|[��=.'ARY��ڟԱ�,��Y���m�X��hM�dw T"�M�K��J��3�i{O�RA�ek��~�����e��P0����6�H�#& (��p�����'5�,v~l�[�uG�P++/3Y��lN3 �hX���)��WgQG:�::;�Y�f�����z;��ڇ�zT�a���� �ɘ���P��:����p�{�X��DC�Ë=����Ǌ��O�ݕ��R�zv�#��u��.ń.�Y��iuG�Z��>�1>3�(J�������/?i��Q����"�A��9)e��}e(�vf�3ϥ�~�K�m=y$��D����t8�OH���rݶ]T(��@��y�<�u� %04Qq�]����s����%� ϼ�id�C=�:��
l⩍:����E���֓y�~�l_��V1=�;0�Qj˷0j��WPʿwqi��m��댿�u1'�I~z���x �<?���w�8�c��5�~lF��p��+M��'�
T����0����e]�ɎV�eT�h���v�{L2�.�t��{<x���Hu��$YP�S����;�l���ɣ 2�P*t�[�����s��d�E�ëW03<
�c`e eITTq�Y���a<�+S\B &5.ۋ���7p��ҏ[c�M�'��-Ѳ�a���`��;۠��w���L�F�]�Cջ�xυc^��h�N�m�2��A�H���3�v��sm�&N���s�S/�@B��$���!5�j�W{;�1����Y^Wo�?br��`d
-�g]le)?��>{_٧�+� e�F꼎'#l0�lg�s�6#W�i�t�i�*�g�l4EѪ&J&�_����1\�420f�ڦ4�䫖Y �κ*����!D�?���%�/�ǕD
t���Γߨ�����Ц�DJ�0ZW+���8/�Á����Z��K��\	�#�Td|׌( ���0ߥ������5����Xso;J���n�L�d"o"k�1�ľ�H����%Bڇ
7z`�{|�u8�&�y8X��ZC��,�s߇��ߟ��U�K�2�<�l?�{W�J:���r�C#�����.���!�8�~!�i�:/l:�d�˜���Q	b��-��e���F��
/�)�7��������p���W���W�AU\�?sf9��y�.�f��Ww	����wG�=Č�z���2*����x ��×˅�%�,���J�Z$��{;^���<KdaR-������L?.A9�b)��4���浻B`�_� � ��Q�@����٭�Q�3m�'3lm/6rhuK��#���֝-�������d�Q^\J�)	ߵ�'6J�� �<n|�u����r�?���5Ƞ�e���0Ê���:׆������U��a_c��=a{�RX_����#+���3Ŏ�}釉�']��K��[�{/����,(Ę��a����ҒƑ����nZ�>�n�y���Խ�E�ig�(�T�fm�
��$K)f�?��[�}�|?�
,R�u:p��
�%O�$TVw$܁C�xR��76�z�*)A�<�1��Űt�D�L�=����p}�̬%��($C�[;�i�Nv�ɖ�T�k_���e�񤳵��_���l-�:N��ޭ�X��Ϸ���I�Z���X����P���D�{�����ľkvƬ�F��PXRXU}z��ZP�/]Fz������&�A ^�8o$s%��^,j�m;���$ ^p+�O�`�8�X��va�ƽ�O�a+pĵ�f�@�b; �0�ėA<��#3�Q*d\���_�jk���V�#W�;lWW`��ōf|u]�X		d�H��cx�D�f,���9�p�T �"D^�Be��0L�}HSRz��c�L��.o)	hZ)��IiCfw�*I�(�������ۏoY\��r7��$R�:d,��o����o1�Q'*���r���J����:,vܳ��$�z/�s�/�4ls��󄓫���� M�oi�9{a.^���"���wkS��8�{G�C.��;��<[����tuucܗb������LiD��� �+��R۵=�]��ЊV�'��Ic�x��=�t�P��4j$��MID�$7��ղ����>�
�-\|�А����D4���8�� d��Uk�#��4��"�?���h���P�����ξ�}�d���~\��t�~��:X�N:����5�J��p9'����|:Q{��r���·�!����nxɀɼ�ҕ���F���+��Hs܊&��V�#���A��-E�^|m�vjf�:v���_��oz6�S��)?�YV�N��wB���}/��8�4�#Ґ%��!|�p4@�}y��NWǪ�c�4�\Ye=]OMIai�m:���~Þd��p���ܺ�_��-��A�<�qʗZv���SU-G��̸ݲxZ���g���"�||p=��RՆ��,(��{����Tȹxf-��D�F%7;���R�@�����W�H6%A�'�X��j����/�Q60���H*@.Q�������0%	J����0mm��Ynu���AV��2|=y�KMޢ���-�g�_�w�D�)�Tڌ1����^3�M���(���3��t���Z�bX*�O�P:�	�f���~�K:�_f�������Ͱ��L��`I�^!/�c�lO:�U[��&53��;�y��������=�Ř9)@��R����r��:X.�D,/i�"��T$KE	�l���R�y��|����`�����$��=1x\����3?~��C᤯������:nfAL�lw8���./�w�r��i�4ZŲo�ۚ�V	���ʰ���5BƩ[�18��,h���Ä����~�#b�ޱ�t'Ș>�KF?�"o���eL��H�����T%�Tgx��'}���fM�2�wqK��#y�x9n�d-y �ANN��C(߀3ZD�����U 6y�9�
}9o�U�NAwt��K�gh�ɣ���0DM<�/��)�w�	�7�&��4��
����O�>v�o��J"I`��Ռ>��ף�nN84� ��t}C�Ō��#��������%�Q�[c��jѼ����xK)~u\(���g7�;͗rVK�Lʫ���x+�$��o�)w2���� Ο��7����-[���J�]�7��IN&:}�.ڙ���xb�'#?���]�_�.�i�ˠ:\o��B�@���ڔ°�Ue�C=�#�ӗT���d�OS?L���vW/4�Yg�~%0�M �K�#���1� �]�e5Y���F�����w��[�vt]�R#w��s�F"Ւ;���+M��#�F�GJ���ڟ-	�}=z�`J �L����pW�Y�� ��>��֕7@>���I�L󄯦<�u�gt���	�O�X�����ٔP���l���/�K;\z�K�<����S�҂7
�+r���x?:+v���WV�S�@t�W�j��>w����#�xU��E9(c���/hEp�u��\5U����������*�QgL(�=2��o]��ǈ�f���q ��,��(QruJ�MP0���Ӎ�����RX����d�����
��o�E�2����_������2�������ߣ��"�V����K
<+$kO�p�n/ �A���J�
�w@q(����	���������0�N!zԛgM��P��o��B��S�����~f�������6!|��?LԢ�tT\���V2���t�	�E�
�>,��QYԦ�M;��@�ѧ��d�v���	I:GJ-�z�d�8���iC��a+�ȟ��Ra5'?���zt>�YQ~����I�b��H���| Շ���[�:(J�ߴ*Ě��f�C�yc%��(�¤����C�ഄ��,!ay�<<be���qbR}��g�9��7���[��2�I�w��Z\;Ǽ�R���3�Hd��݁�G��i�)^�F0�w!���?O���$�n�Yv �v�Y�rr�10�k��w� &���]�yw��|�L^1Y�x�/�1]p��7��} =�ԒS�ҋ��L�7�G���ح%�_�d��y�N�2W���������lD�ad�H��|����O�AE'��Aj���j��1I]6��oL��o�Kt6j=�"'|5�[H4��%v�+�]9�-��%lv��n�m�&҉<����B���lRW�f����8\����{�\�}<$�sC�fxX��l�l"R���o�j%!�������'�Ȱ\p�Y�F�9T�*Ͻ��v����btPAW��W�Mf����1����lٺ�9qީ#|��Ҁ��8�F�E�Ԅ-���hw�I%�Dc��þ(��9��&DO�:�;.X�;5RZt��?X��_8�Y���י��4U��}��5ޠ��E�2��٩�j�{8~��u�FY�XaH��Fc��ï�MB͘�K3L�K{�r���)�X��K�����^�w�Q8R�(��C����n/�x|��;E��y;��2|�$=��Jt��-W�:1�2D����E@ C�=wP�c�$�ߧe�Lɶ\�F�\��P�p��~ Z�ڒ3f�\6���J5n��k�(0Vry��M9u�,1,�h���yw����Cn���&�<�#�$(��#<�4�F�v	$3y����r�Fƥ�~d���e|kR��TDdY�8���ʢ��e^�K͡�mBȏ3����6�wS����L�W�P#�Gމr9�T�ͤ `��Kɔ�wG�Պv[h~]$�T[Yl\WBm�=&;-BX��ZSY��jR�`�3<��Sq�y����K`iN��o�E�h�-2�%�%|
�[1
�4$9,�D�S���#�zC~%�j0�qJ!0��+c?��O�(W���_w@��VyU�7ΰ�3�P�/'_�=_QCp��<ځ��e��#o㖧J��Ȫ�q}N��0��]�g���;j��7S�AMx��k���K"N2�@�l��v5��?H�x����<�*���\F7@-P�J(=�7���3�5ɡ���өL3�K�c���8v6m���d3#ع��}P<�;��)b���|ΌM������)lhB��@���?�'H�Am��Z���2N.�4Z� ̀�{<��*�ZwgmY�M�0.���_6{{�K#��5R�N�[m0��z��k%
S�������!��,�	�v��T�o<E�a�a�eM��?�C C�Wt�Cb5�Q<���@Ѷ�e��+M�]���I��j�ϖ� �˜�G�[�!�G�`�c\ޤ�Ɛ@P.<F�@"��f�#9PM�ʖ-Mn�,_N��.!���Ω�q>�N0���5ş/3XU=�)�ڛd��|���ɒ>n�������o�k0W�i�Oo~눾�W�E�C4�p��1�<m~m�<��W�ǫ�$���c<.�� �@�C�2}\^��2OVq����f\�U/܆EvJD~	*«�L�6���w�Q��v�؂�\34��_B�v�~'�K6��o$0`��ԑƝM�#r�k���6t$2��U"��
,���L7q������<�0���?�����2�Ѷw<j����ꋠ t���&�<�SE���xa��~l����DTA��"`�z?�C��J��$�+��[KQ�1����?�?������o��id���R���?�f�H�9D�N��|��d�i� m�����O{^Y�UUP�^xa�/6��g#dx�(q��k�ݦh��ɕ�l�P�L�<��V���,3^�I�B�3��O(@g�q�U����1��A��vLoE캿{د�pOi�6����}�?J53���۶�㯼Tȋj�2[���go\��&
K ��.ٛr%��D����9^6+�'�����?�2ȴ��#��dP��ڸ���d��ץ>̗Ŋ�]!�ڰ˅L����`������=���7JY�CY5�6�S��{R[�t)�T�R�Xٟ�ﻜ��S�w��BrJ<ѐ=����P� ��Pgo�pw�����H��*,���"��lj��$ɰ#-���E��-U�
����-�1�K��֐uJtM����a��A��O�g�W��b����NT����!�bp���w�c�#X.��)�"��+�
*n�6^b��M�1�} :g������	}��(�}DҧͰ����;.��aZV�U��e�w��L�`�ܿYT#ʓ�X�b�q����.���Q�wb&��|�����ˤ;w�k����}�����ل�[��G����+gpt�+�����-e�P��ߘH]�����F�h��O�[S��BӮ�wa̱�t�zQܥiAU�1Do��t��'n��왣!s,�RS�$V�O�g��?����������c^mD�$�D�q|6��vӐ
��*r�L��4�\����7��ס���Y��sE]���Ք��N�ח֗DVX��@�vp���`?±��O�b��� ��q�p���e3݇2�����D4.j-y��y�f�/��v�s0/8RK�J�Q�nd�y��Ŭϱ�?�?|��{��o:� �%�{�:3Ւ��?%T��UYc���e���Y�5\;[�}���hj��f�t/R�<ީ_?p'+�z���K��!�\@_`u>(���;��><�g��l��]avY׿�t����&�U6n�����Sض�d��#�4�^l$kI�K���+9��B�Z�=���9�Ih���k~���^o�`����N�O�Ic��c��V����:�$�ov�b���͆K8m}Q2�0��r�������/D(��Z���}��W�%�~�ű�矠6)^�Rr��<�5��>{�摵�Р^�4�@���~b'A���B��Ɇ;e�������>x���n-���j0����zjE�N0�������+�HR�,`�r����>H���?Ê�"��y���^cS���ex&ʥ���%����7QdMP�d�}�!I�v��-n��
¯��]K�k���՞{y"�g�����
KOM����fթ��z4w�L��S���xN��~|#dC
LfQa�C���f*M+:Bf�7�~h�&�0!�����&`KH�|�m��Z%�8�$H�ƊM�%K��"JEgƍl(��fT$���n��" ��*�����aK7�n�Yd�����'e�t]c�>}e|S�����Ӝ�&��C�m�d�O��āV)�.�s��<s.ճ�X�<r�hW�n�}�j`�z�i�n��O�$5}���`_�\�;�ZR�q`���:��n;G@�Z����.���ݶ���z)d�|�&�D��`<f��ڰ�_��V)ڵ�#���5�{y�v��`a�^,���e����]�6���6�p�c&<�>�grg9��$=i��_��xL��uEF�
����9{/�*Ίm花S!P�H\)�n�Jk�X/�>_,�\\^'�e�P$a��>�X.nN�aL�GB5��P��	���]��SF�2�]�T�a�ʭ+���,oș��E���}�4%vO_�U�C9[Y친���{������ߥ�z�Ւm!�}#;�d�[��S)ZR�>�����k��S;��,ג"����p���@�aw܅�B���"����g����#x}������ێ��eM�Ֆ��X�F5잌bŃ7E��+�,�v�:Q�&"���tG�h8uJ���)S���>Oy��F�s��Z�>���=�W���?9Z/�2t9�<�[KF���������鸰�U�*%�;�8�>83C��O��b��ru��D|��~?
_dUnV�e�+�W���z�~�R� r���7,��e��K������o�ڌ_|Ka,�����r���ON@�׈�I�}�_g���I����Y����} Y3.��m���K6:�妅nq�sa�UL�{a�;Lć�ֱ����q�+��ˬ��WO���þ�Dכ,��RP���6�)и37�ȸ�G�� �}����n�}8OӋ��<�s�m�$ZF�6ɧ,_% PEc�\ZE�w�ސ�������5:D�����[X�<�#��,�1	c\��HOiK	�K@2�K�������S^���F��8AT�|��L��{�'���hv�G⃾+!���r�^��R!�tOQȀ).��i?ϊIӂϞ��*�v�D;s��N���*��-��P�G����*S���k"�����)���#-nҩ�g�8�e��
��F���bYmg{��iX�a�?�r{���%���xa���W���Em��P����:&o��}�
h�{a�v�]&B����:,����GS9��s���`f���j�ɔ�44�Q�x��5̑X'�8�+t����$�G��K �������Ϋ��P>~~Pcc����z�-ANRn	�J���������zkRHژT�,��v>�9~9�;irv=��bp��o�鵟�0�T_H��}vw�MlZ]NǠH�GfU�;�xq��Zr�tHY��_':�rC�������_��^R���x�J��,�<�L�d�w3�6:�:��������#x��A�2{ѯs�m$��7q)7Y*�y�_�#���.���6g1�/����EQ{���Q����1)�{WY-��n����{k}�n��4@5���p|�=˰����O����p�3~B_a�O�_g.�%�u�86���J`��8���خ�{�q�I���?иzJ���{݇�;����S���׏}�O�����TP�ع�pro{�0�����ԁ�8���6����5
?ƬX��W2�H��>X����� h�@����o�:}D0�h+�P�v{Y8]��ٖU�~s���E2�R~Ⱦp
���'������T15^�^�B2�	�V��	��J%����S-�!omݴ\�,�{b�n��KQ�;N��d�I��?��2�r�~�VKU�s.�fH��W2J���3�
�Ek�s�
�,�]}+R�E��Ґ�wr,*����ΛaO(V�,���wC3�'M�d�Jk���!�/B�_��������v��e�3j�#k��B�_<�h%�-[g����^��y)h�{����
bDn�*r��&���'�.[�}�rp�mN�Q�ybж<E m�
�%c��g�tm���XM�J8{J0}/�DW���=w�:֭#BW �-B���ہ�rz+s�0*@��p�^l ��F[�1Ѭ��D4SyS|�
g����r��]E���o�oeNiT��#m�kG[�\�����k����� gMb�Ϧ	UIk�SfKT8η����!�����SYy����5Ƌ���b�\��v�	]�������4F~���$��@�w���OO_�y\X0�^��ZIj�/�����C��5�.o�<}Yڔ�b�9wI��D�D�=����/�n��V�-�P3����~�;=Lc��l�pFfy,��!���:H����P���L�5m}����+����4lK���c�c�yjV�1���vj�阱�)e��N> �[�	k�
¡NRu���P�z{C�2փܾ#�����2���A�s󖀫%ڙ���U+�)�����aQ��ׂC�0t��H�t�tHw
ҍ�%H#�tw��! ��CIË���;_�u���q�������3�aYע�}x��$�k'~6��x���y��g��
+&�����q4s�'׺���rU�;��ӿ#�t����_��*4�@���@�iYI���w�l�,\`�)�����à���/ k��8�.^R�LR5o��G\������K\ӿY�e:�m�J.�,�ԇ�"��j�=��^ޛ5Xyez�	&'��}��f2EcxǬ�k�������q�8�A��W�fXO�۞�hec���0v��%!�;	���6. ��=BgKkL6k�����T0���L�6������7�k���S>=��0�/@��<3t�'/�q4:��~��)^!�妕S��R3G�D�\qWs���h@ Q�N�%�'F��i U����e�(x��H�ꉽ$LV�:�R(��B�b������L����JSI����}B�4.@�F��L�7�;&�׍��Ÿ�n�l���lEϯ���!�ڈj����Gn��K�M�}���x~?�UBL��Z���X ���������7���X||��f�}} M��l��^l;��!Ӽ�ޓ�X~u
��3b��t��3b<�U@p���G����������%����x(L��]+�G�� �[��/�����Ju�f������*�� �UCh��p�} r��ף��?
<�5ң��Hx��c�� �振L#H��	rkC�����(��:dNܝ�����Kbo��QmN���`������b̐�u�3�bMI���߇�������:�C3>+�v<|����A3^���\���G�/p/�j��ө2b��Ӂ��Qd���j�,u�iIa���� �����,��X�%yA}�ܽ���FX[;��1�$=�2�7b��H�=�M���1�������T��/��Q'�T�xr�W�Z3vQ?��%4�(3�W ��e��� 7�HG>[Gَ�H�1j���v��DO����s�TN y�����(����YоFV�i����j�wJ���K��C�Rwl�0� �DB�Q�cI(����~��B����-<+��(�
#)�$��Io'vi\>Ͳ@����X������pj�Z�Eh	v������ao��O��G���������q�)��3���}����RW��x���P�HtJ_����t�e��:��K�iC^�����B���7��ymq������C��2p�c�I�UiL|����h��n����!��h�Z_{�;�G��y�H�[qy�oǔH8�=�[�]�5�+|&4�}|� ��f�.o��iB�@ʶ;%��RG�{��A��Q�W��1�g�$��h��큭��[B���T�� A&�jc�}38WZ^�� �~�� �W�"<5�eۙ�TH:x��j�A2��b\��2���p��n^"s�IX����8/x�4���yE�a��>z��}q����l��jn~�j�� 1p!�D������1G��̶�v?�3$N�O"�!(��f�w�!�G����}�ة�����m܏��.1�V
qͰ5�.�y!_'���f����pa��3�T]�?c�?�?k8��Tb��l�.������
3����3��g쐂OF���rU�,%�P��="9~����#�Ԓ�0$��A�T��"��_�Mɝ���\�85�;�m{6��|مN����=/'�72�/b�B;l���3?a��1���ey]Խ��~ �Z�,�1EA������܈)$�s)�;^*�H;�X�r#�m��Iv#H�X]WߊE�)��L����jў oȈ�^�OF
�*�T��=$�	��Nޱ�#o�E�
����3εh�l�S�z��v�>�}	����r-MQ��Eo�w�(�o��T�[k|%��};2=��uЂj:���^�{�����w$�#�����\Y)� �����
�j����#�C���k����0�GBd�Ҥ@�5jV�(������o�Ϲ�=*����v>����i(Ʀt�2,� ��D�v ���p>��w% �5h�:c��*R0�C���Y?@p���ܣ�I��+R�d�a��㢪���3��G�}����?d��.4t�$�>��%z��2�vy�q�{���Y5m���vh���{p��ά��+��I�����K�/sN�-�?��{�+��EGJ��ϧ��[7�m�ѱѭJ�lh4
�/�R��޷@F�r�6�7،�kk�]�[B#HL��7M_c��t����Rw�
�IT@�x4/t�^Eё{}f=�A P�h;����n��5����f�W�s��TW�)�!r�ų	.���f(�4+�mi�d���P��7�A3�JKO �O§ʕ$�8�7S/�`�~(�z���pm�����L=�	��6�BёNrاx~�:d]l]<���i����&gfC8{�Ƌk���ۙ�̂ފr"��3u�p{C���1`��KcEW6\j%M�usa��1Y�J�g:�5o�uQ�=��H���-�ϱj�Y�>_L}fɂk��ئb����}h����mGc��I0��&�G�銖n�us~Z��'m��ԑ�z�Q����k�6'������ݮ��ý��U佼Oꆢ��yŒ!�'�����.��ɐ鏟�J��N�G�	���W�ξ��4�!�|�:�kM�C�y�V�$7�[��0�$�_T8SO�3J+n�϶�-�n�;�_}+y�w�`ʏR�ۅ�5�o�"!�xO3��.����Z�҆���9����aB�ѳX�����:<���Ұ~�w�{&Ku��R߄�~��7T�Pv&%�M:���%����zTcB�;�_�B`s������S}��g}�!���-fG1������X���0k�*����o�aO�.�y֦�3h&h��orߠ6;H�a�ܔ|Yn��p6Jzr�=�,�B�M��w�(�I�'�9r�ۼ�X|l�k��&���<G�����Ƿ�]��4�T�<*�h��qJ��®V�F#&ȍ�F{��۶6G�(�7&��| ~�*��A���[��S{��JJ�,���H�rJ�]�M>���RW\b�s
� WHa9�b"�G}��Q����é�u�М�I�;MA��=���D�o�۝�$;��Acs� �>tq�vɦ��>��(��B��3����Y�
'�S�͘C�=�/�{2�tϗPo6;l
x���]���E�E�9T_O�Zl����9�ڡ����G�H�m��<��ə�S�6jH籤_�6'P`X|�`�<>�V?��TΎ������t1�t �$�NA��i헙���Ӛg�Q����� ��Ye;U���j}
|�&>���Kt��\���z플������Š�;"�6&5�V�B��g#����_�$j�ID�p~0�І�
Rp��|�|�2Y�+'�Z ���ZKk����3I�������?���f�/W���,㫷�1V�Aލx0-[���~QN�����˱z�N�F҂N�1��T��34�y�� Y�<�/7�����m�*B|>77�_�5�T��Ｚ9{\�a6�w;��{�܍*�%<{�B7�7���I�pjH<��ZW�k�n��^�ɞNd#���B_n���b
mŉ]{�_1z4A��0��vPr��0�6��ښܨ��=��D�w�T�x��qo�\R�>쵰��	R����������j`�ZHfC�F(��s�E
�@ J�#�����6v̽���VWj�-b��� ��4��|�d�_��שH��IN(�ޝ%E�ɤ���Y������h�=�>�����pJF ��gT�M1 %�ک��3�wj�UE�4��8�F��_S�xWC���?:�x�����~y�_V�k�ҷ��FI��gBB$�V�ʔ��k1a�=Vk4��+����.$��+���s�M������b�b�������'��4�����q0ԍ��a@�.ͼ#'Rx��Ug�PI%&��M���NY����S�\�=q�(�����u ����2 �PG�?L�vBM�G)nJ*�*X7\������4%�c��[���<�~#r'�}��命�'i>jJ����5��	��CB5E���GA���RA�DҳN��8&h�f��.�eEm#D�C��ߎ]���ϟ�C� Ͳ�����}���?�����AΤ
��D���#p��԰�����{�׼q��0$�o3�7��c�D�N�\�v91�RR�����5A�N͆�ެ��O���;'jm̧�
�ճp%�Gh�/��aX � ����_X�G]�,j��˙���Itc�s#m=�s�NDsnMY�1 ڟx�^��9������۝]���0[+����Q�V�_h�O���懃�:���f�O�7Ĵ�d]R�u�i� S���W��I!�t7���$��E1�IZ���qv�XN�-'x�[5��|�n5��-:��3�J_z�cQ�t��� E �"�
����M
#���}K�{'w*i���7o���ajZX�.�=��ݖ�J,롊��E��Jv���+N��*��O$"�,���Trc�;�A+B��� ���!�����,G���~`��U�`ĸ�/�������n�NԿ�EPK����Z�o�L%͠�����N߀Z�)M���EM���x��6��o<���	$�%G�M��`K�`;���퀗�=7	��<��,M��U/_�@����kq���x��"|:E�G��E�[��;��Ҧ.%�@R�^b�\[{�y���k+�D��H|�]Ŵj(s&8�24jEC���-M��a��阖�HV�O-a�I��Z~_�{G��M�VX��I�O�ŇΥjV��d�U5i۞W�E��?���"���b��'��vی��������֎|[CT'B�;�Q�vј�ke���%q�Th�̇���y��b	�͝7ƛ�W�}�E@)XG���^�h�h	=��8&�t��0���u���� ���oS*��t5h�S[�*�Αw��N��EOn�`?�x�
g�Eu��3��L?%��J�T;C�oM��&��Г��-�p�q��%[ց��k�=	�7ZʼI�]m���!t�Af��d��9_���*ȉ .��t����pkCrh�)���*y�7��U�:��<�]�*�&�y��P�@�w�rK��kǂPJ�(�g����N��+����`,�ԾKL�K[��%�2jZ�߾[/J]`*�l*���z!�ê�&�,��P���E9��.á��Η�d�KO`bhܹ���F�S@�<Џfp4����������?�<����g�^��`C�̨�;�ͷ�RAB��7}X�I�.���t�^�a�<����q!R��w���A�}�Mw7����n/-槝f4�
a�Vp�N=����+&#:�\�x�<0�V�H+��2��VDϟ.�;�iǧK��ly�tE�w��6q'��i�-�g��g#{��o��؅Ј/��Ǧ�k����G"L�R9�-��Z)���ek��}y��q��w�f���Dy��z����n�f�0S��tқ�Q<�3TC���I�&W��.>mG���� �\����&BП7��ήx&f���PrP�R��������a�m,�>xњ�Q���s��,xe_��"�3�t���_�c���.<�E#��7uM�O�X���vų^g��F�Nɒ/�W�"��:����7��BR�ZI'�3����Z}��5L� ��+�!�Ӣ�,�2N�o؉]�#Ȥ�U)�m|:9攻��L9����_�ft_78
Vȴ��[�x�4���4��F���n.$d>+�����Y�����b�]�h-�ǽ_%����]�UL��.>3�Q'K0��zº�T��J5�&K"Q|V�h����S�7���U{��	��խs\�&y���3�-G/hJ���������M��3���ӧ~#�
 ����3չ�?訴��!¬8K�j�s���1����C:��<�+Ў����o2%�J�����7|;�:�>,Z`mJ*�A�j���b�'��5P�"�;�~��$�$:?I��rB�kv�����^G�����D^K!�jN�=�zC�^��SG��~�;i�`p6�M3�[�G���/�Km�SF����"�+4r�g����Aj�#p�OX��Yurt��/��>�D��-��y�����.l1�T������2���
��̒@�kP~�T��»k}�㿻���?���C�9b���?Q� 8�Ϭ=��H���)���;p��2al�Td�!e!�塨U�'�gF���[�ш�֧��論�l>!8	�TZN���u��Y��/;q8`}q��r�b�̆��U@����/($3�� �������|Twudf�Ľ��+�Km�8|�
�P4�)U[�
O5=���R�P�vS�^}k�*�@�\<���d�ϯ
#����~d���z�=���mz3��p�HL�`줌��n	�՜��T�tՁ��a5=X�ru���̲�����olɖ"C����=C�,*�c5-
����rDS5�z1!��~%t���%�|$O^	"jl�
�*�����7
���r���;��˃R�$�z�,..���<�ܡYl��6c�K�~ܔ�u���u|)܎`��i&�#����]R�`ƚ?������J�m����P�� ���!"hPD�	ه�5�4����F�B���q��{�Cr��dbl~�Ľ�����C�jF�W���}~3�d���QSyKG��6�(��D@$�B:�7����{�"S>�V�4h�Ic�8J��`�N8ng�}��к��0�c��T	�[-�d���m:����X���y��&��ʓf�B��	�������H�vYxXD2�y��s�.�gk��9EO� �9� R_��%/����m������RP1)i��K�Uã|�4����"��!oP��1%�S�V�R� ߬������{Y�����@wTa�����31���hK����Z�*���,���7�Pj
���z���2�`�S��}��*%�sxl�]�8�{��Ci3'��d*�S����Ny����o�~`Y���y�vjT�DR!�c�j�{�>���gw Z��F9�C�˘�`�xZh�"�����-=R����Hʬ���,X$qmܨVh)�'�k�7�,H	A�qV!K���\qv���ʓ���U������:�W���[>��G��q�I��vP68���nu$y�� F(��MW5��m;3��J<�O���=�'���_-�Ɋa�/"��Ĩ�7/��I��y�)�&��Q����jS��JW�%.~�\��̾�L=�u�g�"�u4�r�!syz�A��f>�Ԭj�32z8��fɘa�x��v݁,�?�ǐ��cN��%�n����=>p��?��88<)EAw9����4 `�<2��?�����o8�{�����ô�O�z�Z���;�n�~u�av�~ED���˿�wɘB�83݉�r$���yV��6�z	w��C���=+hOQܫ��\xT!�*�G/)G	���&y���F�B�k�a;D�Gf��'����j���mo��Ɵ[�(�vu��T�����E��[P�.xM�&(��t蟠�zc����De��P 2	|*�8OmX��y�"➄�z�����EA���y>�1�*e`����<��[��ϛ�er�!���pV_C߾�z<z|rR�L��|���&)��X�| Fvu@-9(A/V�������m�������bQ����Eý��A�l
{��s���#ޛ���ن�x]�P��u� �0�7��\��Fq��ꡅ�&!��w�lk�v�`�\i�bՐ��+N�ow� -2
7K���R�T.D�(L,Ud�j����ƥ��A~����uu���R���0�$d<�0�E8�:
F���9�}𗭰�����$��SD�9ӆլ����� `z�D�����]e9E��M�h=U|�HdJ!��:�#���㇜8-�<�`�F�\DQЎ���<�X �Ar���똡�n�b�����t-�\��
�j�)6yS_�/����s�>k6(SB��G���Ie`��a�ћ�.�� �=�t��OL�
FNl�rӎ̠8���51�9�o&�K�K���m?� ���>�{9��Wm��4�tV �D��
m�$�3�&�N��Q4��a�����+[k���"���e�����JQo��v�Ⱥ�wX�n�tk��W�Ź��SQ�7���n2�z��8��q���w��RL�6d>�-�����!���ۧzv1��K/�Ds�Y!e
)�5+�r�aU��[$�P-9�_����&�M>�H6j��c�YE ;7s2�ѭ������N���K��n����#33�pF�q�N�f�c�U���#U~,ѭ�� C�8���%��Wq�H��w�q�5A�p����,���G�R�Q�FB�� �z.׬W�D��+A����P��ǳ�=��H��= ���i�;e/|=3p���P�%��{n�4Z�di���[�0h�5;�
���S��ٕ�z�"�L�������UwFbV�A=Mf���qEt� &:�:�k~
��.�L�#�-�9���
țI��U3�k����]щ0k&i�V{��W�=^S�W��{��\��J]1C���t=O�\�����On:11�[뜒G���ihI#������>�mA�]췲�l�__}�z�x�+���R�;���Bˍh������C�CD�����R��ϩ����Ď�E�n��4�r��Lw�r��Ė�!�y&�:�����Q~���L�H迉�h��߅t���^�f�P�$3D*�$j����KpR��h��|Lk�Y� o���+U ��P׃l:$SP�Z��P�wt�[��DY��(�5Aٜ	�mg2*��|��M(y�@�W�^1-�ޢ�o;����2���7�r�Mgl6�v$=��%a 3yw��\obQ��+
�DR*���t,:sj0&D�M����u�Z�6��9�T�$U�VO��fY?�~�|F�K6Ìiͥ,q�L4g����J��d%�������3����nT��͈�1_������zpҧC�I��$ q.�S ��w�f홵JF����j�����9�)�T��ط^!�e�T^�E0�E���ط��dN�54��j��(�g��� 8�H��k� �_��d�$��69�K�G9�9_���;	��V�rhK�+}���P�?�U&���:�>�ܿ��g�B�����9w���*��1����$�ȝ~7�����(�@1��<�V�Q�N�FXݴn�d߮�B�+M��6I����ɡ���B�:6�Z {��񳢿����3<�K�$.���%KwqKɥ_�g�9)�	����zQ�Gk����l}b�`ץ��L��Ҡ��ަ
�9n��])��F{����W���2\�s���J�r�@��w�3�QMF���mH(�L�VXH�]b�Y %��G6��}�'�TF���e|�T�+@����Tlp���"P�I����uxh�`&�5�>�z��,�V���q[��y�tHP#Z� B�J�{VWr�1�m��v��)�.0���ۧ7�s�-�Q�G3��;��R���鯝f���_��z�U�����:��洧//��v�(~�5�� )�=2<�:�La�&Wp������c��7���f�Ng���G�$��)Pf8��8;k����M�N,��"w�#T�}��9�W�v�����S ���GP$��Z�;|��� �L" /��ދ_�/̝>�"�I���Z~���Z�]Z�[>�įf�/%ˋ�}��[��żbM�,�}�a0����X�����La����"x��C�Ok��-.����X��0c�J����&�c�a\��'�Z̖1M��/�f�������j���o��;��c�
K.���Jesb������:+�?3�{�����*�*I�����8���w��Nogyӯj���Qv���߲8���Qrj^u:�9S�>�f�M.�̵�r�!���O���g�g�b��>j�+�-3�VD�յ=�8t��ÏTo�=�_i����,�f{V���@����4��K�1}Q�.�/c����$UB����+E����VP1��q�r�o��N �GM�^ۿ&�P�K�,7o�-�,�C�k�G��O�t����]q�kkS���1V � 19�_9�6>�D���ԁ�q�`����D7$/Q��q$&���M@��sW��&9����<^�"E�h����g�����E�������m�a(Gm��s�����l�C�o����Kܝ'2}�B����Dx��m1s�V�FOE����5��I�O��U��I�}n����xOUR�KԞ����zk�q� ;P�0��@����U��y��v�11}:�}�����+���2����W�C kJ����u�r������]-��@YWp%8д�Tj�����/'�����'���������
'��Tq�����EW��ĖFC�z�����#~*Y' �m�~�B�u�t9�t��,l���^�ڱ������vov�M���_��&/�F��L���z�f���F>��������_9ٍQ��\����_�ۈ�Z٬0?݆YƧ��F�Yb��O��)�pw�uX��r�(�#����9]LF��Q�Q��n��Ms����>4��;��<K$rQW����$���RD�%{$�Wݫ'ϰl��<����q`m��U"��/�O���/�c�#�?N�rQ9��(cnƕ��cgd��#%*Up�k��m	s��uQ�)~u��v�wY�y
�Bu!�aɓ.�>w��H�	��wYD:��8�b�M�ɶZ�SV%���[³ l���㣷�B�ЁɼΗ�@�u�V��Czb��'�\K�_��g��O"�.�vM�.��3#�V6�,��Ľ��� ����\¯��R巖�B�S�'��O>X�����]��H�!m��DM�ju�R
������_ܞ��	JP���������t-�g�@kocozRVt��'S �����k�2�g�~1$QNlZG bLo���y�s�;ȹw��6�h3�EP��s̯��;�f�Po�f�����$y-��%�W�y2�B���[ZZ���:ѕ	7ͯ�	����{�r�)/q7��/�0����t�$_�O?d�D���Q��f'4��5�a�Dٯ�t\`�?9�bi�]�B�\�lƶ���y�[uB����e�~�8.+"��{yP�ݷ������k���﻾u��S��N���Qp��?�d����A�[h��ֹ.:^L�"������nz<>�B�8�<����$��V��N@��y�+��]fz���D#��f���V(g5�2����^�GP�`
 ��=�x�������2�9n�ө��뻵�"N��m�U�		��Ml���XG����O"-�����29(���g�{l�Q?��Ÿ\�}�������m�;�Bc�ngM�No�$����6��	�6a�H1���Ծ^�7��䈚?t�Q*e������������؋<�UTW�C�$E締�Z{u���m�HǊ����&�E7E��I��X����#�l����Z�f�k؜@N$W��[��9er#�)�Ց��}̕�p������i)5�=g��h��6n�
�9�����;;q�G��s���*п��I�@����=�yG���dY�����h����x�!�{W����x'`��+�v2k�=�Du�?��QE��(u�������L>�L�[�.`���H�T�Û�X��j~��ǈq�O�K�g����.PtD�w\���b�<��
c��:��� rި��Ve[ڮM�����!���T˻��m�5m\ěZY
uJ�[gy^	����(�Y��H�"`|s������WN�uI�Ǚ��t&���������(�UR�@��˺��$Z����t��d����3�1r&)e���'�a�BTi�4��`K��<(�l��)1D��O�8�����Q0C��f�3�l������>�Ew2G׺����t�p�Y����G��%����0�Rv'֨��(H.]�.�3l<{�/^T�ȋ�с��<a�1���ϋ ��<]��l�6��b�.�ɢ���;ɏ�����Jv.�dLDM&I}����nIy]:T�`��ѧ��S�,��jH@%Ϝc�5��!a	-��r�i�'��+6��0s�xxT�I��x���aL���Ma��;f���2ؓڃr�|��ujP�q�Q����p6g����.]�o�I1�����-���t�ݕ[U�fF%m�;挧�������G�*C���\�{smk]T�ʱ�c�w�"�3�����'�#������d���P�+ѝ�O�w�]�vI%�@�\�6�s8ˉ������,�ӎO4I�b�>n©0޻�&z�`#��O�Z2�O���HJ]�"�][���5�ȴ�D�E\/Q���������t1X��� P"�_v�}�u���J�i�93w��zƅZb5�L���Ծ��0��h��F��ܥ��$�V��_ ���x�����nW��ʾ	�_��������F�s��6��r��wY��1��|�bEJ�g�t����4�iL��M|�Jp|R���:�t1�O�5�t���Q���"�������Nְ]�C�窅e����|Q���(�)'cFo���vo)��6�!q�/�}f &@�g�gM����a<K�)�a�H�TSV��ʤ+f����V�!��<��|d�^�_є>#l�z�8^|[�a�m-.�_L7Uk��a;��Z[	��4ڑ>Jp|6`='(l�*�MƴC�X�Se�MX��� ��T���ACr\��'ecJ2b�����ydl�܊v��.Q`
������`�X����8v|3�&����-�\7�XN���1A|���g���ȁ��$˳.�����j�'�㰪����]���U�<�}`���D��ϰU�:��ֆ�ִ5�j�ˆI�[Ӭ7?ڱ���XB1��*��bl����3K}����묆���T����a�gL�BR�a���ɖV��O3Ҩ;��O	�c�t�-R���5z3�j�WVF9��a'/�id"G�b$u��e���R�ؚܸP�������hNC8�n��tU���1��<5j�(���0ߙ��,I�2i	�����:Y	�ooUh�z�c�xn�:L�)�)�NY[��1�}�eL�b0/o9�I�R��o�-�'���ֿ��Ź�  �<q}�r�C�A9�������p�ח�syX�-#�p��$���	vL�P�^Al������{>q����~��Xv9n)���:9���kri ��a��^t u�j	���)ez�e�hP��A�Z�?kG ƾ"G���۲m4�;!���}8�
�@�]<�e*��\��m�k���`7H��x�º�_s<�
�+����x�p{�A�x=q%�Ҷp���wx.�1�|�b��G�._�P.W��c#<2f�hkY`����3��i��79k/)�cD����Q���4�7Lh1��0�e���8�U�xVe��j��1��W�eL\XM�6.P�w�y�P���B�Roމڙ<ş��bh���}�,�仄0և�Q��3�0U�*��~��1��#t.�3��F̉^��,��(����L�_���t(g
�b�J@{f�]6�D5����ޯ������tɨ%�&�2�w04C98���񪣕	"�f��n8J>�9hM8�Iih8��_����j3Ֆ��x��f���/t�E�K�^mް��^ݨ
qS#�ɯ�2NrU<f�H
�k}������������_F+��/���f��$1G�o�BBQ���:x�7Ȑyk�%�r縷R+��jGAׅ�B����ij��/�ԣ�`��4��|�X8>^�_A�Ц��;�6n;�Jv>�-���@�����DЌ6٪N����m���Q%lmC�瘏�?���R�O��)9`�+�8+�����s+\�J���隔��,����D�#hu�d^T<���̎�����T��rƮ�W�Y�?I�� P }��&I|?2��Rj F�8Y����g7VXx��'�q%�g��Lj��L�ݐhp#/Gn�� ��b\M{O{!ĬJ1���ɫN<Nz �Y�a�}3��8ȹv�e\�oP1
�c������w3��>I"�3f8g�OJ��`C�B�atvҌA�a�A{��'�?
-�n�E^�ND��¸���)���3�z�E|+ei�y��*��u���&K���þo-�|����$h�'��� ǘ�r!.y��8Z�X�&�8Vvs��u��E���Up���� RvȆô*��4>'d��.����.�4��u�b�T�JO����Qf�>�l欥�D������&��K#x$Fbb  NỡW����gF�d���«h�U���0�1,�	�s��;A��2  l���HA߳�P퇭��&ڎxA�������F��8�8�F{�&�{�h%�ڪ�N�vO:)q�Z����]�NE�����$u��Lҏ8�=U��I�bq���l4<�~W�X*-�I� �|�"b¼�K��Pf�嶍<)���4�H-�"��1�j���I�l���t���a�����u��<���:r:�j$4�7F��t��)/[����X�^�=EX:ϺmJ�M���'t@�X�"ɓ�I*�QEA�?�����\;	��h���y���I"���|��U�Wȉ�v�^?d������*�<g�Cx��F�X�H�rz�C�ko���/%m���O�m��wH���Z�@h�l�.���͜9�~���d&��>�\���JCS��*�'Y
�Pn�S׉6�ć�PT�V:&z�l���?���K��I�EJ�:i?i:����C����Y	`JnXO��V��Y�g�Eo^��<Q�_)eN��jk����U�9��gY�k�(� �m���V���]h��p�F��T� _�}@���6�#<���z����4���'�$m��	���4�sOO��ȴ�a�դ
z��٪?���6��F������� {��t��[�`�ӵ*��22S������(��D���(%��=����h+�;NX�"�[<��}@H�xCҿ��!䟣�_^I��;�	������ΦST�~��jǦ���6?�Қ{�2h� k$=c��^ע�]=r����|Ɏ��J�p�ة��A��gJ�0����cu�TvW#䵦]����-k�T���e������8[Z_^[��_Jn�:1���Q4mZ�#@�%Ͻ�4����Bp�cjD1ujzw�3)���CJ��֬g���8�)п��ܜ���o��٤�) 
c�!���+��Lê�4�}����}��ߴ�O�K�_�׏�Z`��d�.��m4H�%����CT%_�7j�μ�^���MO�Ī.���%��=�*1@w#f]I5P��`f~_�}(��T4���&#�AR�]peH��t��e��:��UŚ}'�P��x�ioȸ�z0ԭ2Ĕ���>��ȗ90�,��n;5̐�
��kqP��.���!�6��#���!z��%���H��ERз�-��|GQ�d��2��9_N�	h�%q�1
덖TM�9�W���mH�W�Y���l�ǽH~r�r�
n=QH��k�XB:��?�y���K�����JEk-{�.�ߙD&_�k��e�SU�&��C�lD�="��#��2��jh�˛�;��9	�xs�6m�7z�ɴM�� �6�����{����s6G��w\�7�JU��%�]T���U辔��qjL�y]��:_�J��hOt�y��<�n7c�7��H�՛���f���k�وbSB� �8�d�Z�11&7R^��&K�0�!�����ҁ�[5�ݻ���ku����P �D�d连���m��;��L�5�)k:pQ��5]��+�y�	ϡ[�s!�Okh���R'��,�=bE��HCG�]*�����b��EI�M��*�~t���*_fϵ�����l�P�ݦW�����[�ʢx���1�� @�?�@��M\���zM��s��a[ikD�L�'}�ջ@�B?lJ���Cf��U�������`� 9c���D��f��4�(>�8��/!<nĘ	V�t~}����rj��M���M��;/�VV��A�o�����xڰ{��'n�n��v��ͥV��=��ُ= ny�HB��jh`�c�6�w�y�tw�����$�;�c�_Ԋ�w�p�E�*����F���C穐�U�*j� ͥ<s���-xv����
���X�Bqw=���w-Z��)�vpw砥��ÁŊ�Kqw��}c�����9�5�#I�6� m�^W�P�knZF9�*���/`���,��˿D@R=�U�m���ϓ�ɬ��B�a1�S�{�~+��a�"Q���&�Aז���*.���JK����ؽ��@�P��Ș���b[�S�/������SJ��7npr|ػCb8�4@4d��gd�N��zRkR9������U������ekҡ�չ�P��8���TIwZ���mL�*��m;�V���i"�e[լ���pM�_�,�IA�ɫcE�w�EuX0:�'�@?@:_����������&��X�ֺy�ٯXS���F�)r�V�pF��sQq�}���NMr����_�,�	�g!<��&C�zVbS�N�&�[�o�?0J
e���-Vi!LF{'\D W��3|5���"�����-#A�s"R���4�F����'>���l�����F3z"Pgsڶ٨�������f<�AB�.���Y5��#z3vr��8�����V�
}Mh�Չ5(�1�{�FFEdm}hY� �x�B(�E�v�L�xK��A����[t���K�"��F�z]>����L�����~��;+{�E��<�Jj��|����w�}���Ԋj1�� g&�f�+����wM�bEJ��B�	i������x���o]�3X���5쯥۰�z[c�=�8��&�3X�u�oo��!w&��/��f��d�Y~�qT�uM��%4dfݳ�ɪB��7�o��_��1�6d���[�0�A�i*�ˮ>�+B��:bu���yceãOi�fP��z�߬p��TK�LNBH��g�}3��&�9;��S����k��{�l��a��� ����VT���f��$a3��Og��ƽ�_t�?����W���ƪ|O4d��I��j�Sm�P��L�5��G��>Q��`+�MvO�v<�����hq|�r%�o�⡦g�|G9���D(q�d�O.��'=&�(�:ڳ������L�<���Ìu�tw]��_���oe�F�W;X;��qD��i9�Y<��I�TcU@��O(�7��IU���%Mu��?(�����&64V@��"SeB���j�>�2E	[X�Cb�2�����E25��u������0p�g0½Λ7��jj%i0V�J��|�w��8S��)p/������{"s+���+QN/X.��+������w{��=�w����j	V����#��"��=��%�I��n(ߟ��͎{1Wi�eG�z܈��C
�t���/�`
E����r�[d�PΘJܜ�'����9�EWE�#6�VB�r�"��7���k[��
��ru�#���sҶ��v�w�cpE��MB�-U��d�8��~p2od�>�?���7��+�"�� ��s*��byެȧ��9!-z�+M���i��4Hvr`�+��E��'��a�EOH=!�"�x���J��X��iO���OK�&{9Ix�ն?���J� a�����[�����~���q��D����8O�ó��w[&I�H����6���{'2<��[S� ��R��	A�6)��LY�l���>B��5;�\[�e�i�� ��!EF]�v�e�z��P�a~IT��O�A�o�H�L舤O����ոt�{G*�e3p��ڱtN�&�V�"{�e�t%?��1�.�Q<���]�}�z�L�E�j��O������vUY�x<�G̡���-S��� z�+��ui��ۈ5k�^����zq�PM}c=���ܷ��7!X��`��t'��n���kȥ<]=py��*��&�9�"�}���3�[ˢ�M6�Я^�z%�F��e��3�
��-?Qc�۠8�@���qϠ�K�S����:L#��rB�*g��~��ڳ�߾T�M�3~�>����k�j�^bR���M��k�	�+�Jh����̫��o,��^4<�3����Ff�w�v*�Ga�i3�-��rr�W�Ѝq�3GR0��R<$�ԙ�Ti6���bIݸ��w��u�M#<?Gnk����q�m������6=��58��`�Aza�	~�bkB�d4R(w�ԁZa�B2Y�hC���K��OxFjs
	�i�@5�W��]~y;�e.s
d�ׅs�3�IqlJ�I?$6"�+U"1eZ�Az>%���A�{۳Q���
�?�ϒ��{� 4Q4�Ŧ.>�/'�7]T)2�;?~���a}i»PGG-I�-ɘ�>���j����3Q�%���I�?
�Q��Ĉw����|�
�Дa�O�������������#��U
�D�sAy	�rSI͋��[ǐW��>�B3@;Sk�v��ұ��,tq�i��q�������4�!�����Z����,�s�I���+���*
��$�\�N���A��^B��
K��\����� ������z4�}n�闵�F0
E���#Sʺ�4����R& �rα9@�Ԉ��/�Z�;�]DU��#�����R�oړ����'4Zp�0��4i8��O"Ս�X�8*WO����,4<E��J�����2K�ͲvKM�Qh�S���\<�m)�h���M��|`0ѕ�_ӸJN`w���x�y�2�����
IN��{�h�A��+��O�N��^�X��;�{�/�/�o��M�l6h5�^�~Mc��Z7ey�"N�1���8��y��%[��������,��ղS��Lj���R�t�<R7 S���s�/�h��_C�y�_�*C�	e�}�^ �;\���X��Æ��aBf��ц��Z������b����*A	mP	T�"j�x"�)*�1�#�6��oa�^��!�z���a�)7g��GA$;�	@z=�/��P���jbW#s�]���6�&A6l�WJ������t=%�6a��L� y�Q�����mOGi��JP�d�6�hEy���p+��|a�Gtj ֬J�_�6p� �*Y���<�M����b3�6��o���oa�L��V��3��4L�0e����~W�'4R��x�b��Pe��U>2�z#�Uv;ٌ��액�½��!|��0���\\�]�� �t�LL��y]
}���G[���K�*=�g�kC����0�D�7:���?2�4���t�����5�/}�yG����崘��G��8#`<hy�g"G�LD����7��(o������*�ec��VL�h��T����<��5�H��r�4��ޡ!��Pcgd�5}bt�����m�/���4�;�m�q2�+]+Ƙ%�顔�F����l��~:)�	p����6Ż�:j�MtŐ�Q���(���Pl�!�mv�����'c
� ��G��V[Pj�wp]�m|��P=�Ά���$f�G�ɫ ��
�C)��-R����.�����M��
���a�,��o��r���$a���N�1��*L�h+�y.�hP4`�osܑ ����7��l�^�Gf�����*��+>(��P��fI�l��QҒڴ";%�H1�L0G�(��f%e�'��
�7��%�7��c�#Qs6���M�%:�v�C��;���s��%ê�EB�rb��<��T7������.wϊ4�ြν7�z��K��G���L��l<�gj:`T��U�`�P?�R��*/sۆ�c�E�y�r�,@\a%� O�tlR�K=��޼�7�'4�~d�*�H]>b���1P�%a��T�e*�HyeF��Er5��p�"��g��1�'��&x���K�%�9�A=�>\�9����
���̊Y�6��>P�GE�&s�!�rQ����j�R�M���
�acG%�| N<*�E�r�P�/��3��B��;mL�t���8�tD�D��G�`K_z�4��-݌�H;�M�ŉ��oы�en�]<ߟk5`���}J���\e�*ɡ�M�}�n���jSCWy,�B�{����j��1<��{6�>}��I�%�VC�c�4�Ӝ�kF*�5�
泔j�E���|p%�#2g�m���C�5��,�	��H�A]RyhW����s*�����b�A?�ݏ�I�f{4��	5(�9��=�P�lNl��3���hP(�|���S�@�o�+�^r7��[��]�,�tMNQ�&~؜�:�p4���=��"�;�+�=a|݃���p�P���><Q�Q؝��%�#�{�O��}����)�Ǿ,Ș!U�C��oe�&�_�-F	�*�r;u�7��x<Uu��L6� D�>� �}��4����ء�ܧ=�+(���Nl6:����Ai݄WkD���6 ##��8�L����a�l)��M}���#Vtb
Up��S��s���רnz���r՝]{�a�f���7J!#�f�Q�6?Q�S}�*��-WG��ڄ��1�%a�(�����s��m[q�f���B����Χ�9�}G2>/���*O6̄+� ܩ�[:�z�U>���)l��"6�CLK/~=��F�t�NU�4��,w�O5�W��DG�f��U4��.Z�A����TU��_1Y�����?�N�rut�iwO5?Jh'[���YJ�#%}�$l��Lƞ����ȕu�T�x�56Qض_���֘d���	� <p������o(�l�7=����q�d�f�b�=��L��W���v��9aMd��?�F5&��{�D��1��P��V;���i��H���x��	��	�ݢ@#��G������?��;s���{�~;C�N�ՎE���
��,��<d�R)n�˺�[�F�i$�W�Qg8�`����R����� �ר��~80W�)5�?�Y'?�pxF�c��E�ڭUYI�����!�h��íeVA���_kۻ�[A�8â;poX M��M���������oSK/�N�?t�-�W�f%�*)�qN��)4�g�Q���5MJҪ��aċ8C֤�;F�oj��� �����o� G��YW,��ge�8]���k�J��/�6Pq����^�WE�<����4���|^qXW�C7,WꗗA���aD�G�w��c��e��G#� 9���;Ov#x��T_����"�[��QCR!��v_�N䢍�rF/��b_�sIT�����4�iϜC�?��dwI��������	����)~������~��$���Uï���L�y%)
!��Fj
��Q}�Ԉ|& �M���*�HG�M�)��	��G�����%|P���ѫg~$��D#� �e�V��s�n1����g���v��ܟ?��kuR��viw%�*7NV���{.v���V=ߨ�fQ옦�`*�H޲;=���W�����7��隦~V���|��H2��ؕ��9<��H�A�mr8S���`��d���v�ĕW�>3��j��G���+�+zoLz�?#�������cx��M��K�oo<�=@�Ϻ�9g"}��S�sjV����/��������[�������R*4ͦ�"\I4�|c�P@��dp �ֻn�������j�}/\\⳩�� 2����Ő�a�Բ�w����ۻ�	��!hV���2�N���ܯ���vI�*��nX�9��EKU;�s_��l3�Aį�\֔����/��	��V
�����mM��뢂���pm�^N�3/LN.+��{!�z�.�p�[t~��>���rM�4/�Aԅս��F�zY)-�LX��8iJr�}R/��}n���&Y�\&}{U|�3��2=���<iwNEwM-���W1�07���0����e������G�(&C����J���xV~�u�竭A��Nyg�[�G��l=}�=RS��,I��-z�~��rqt~#1�Zɜ!���̧�;�Ă�Sj�����'ʋg\2�9<>�J�]���P��ެ�hIU'�c�K��m�����9�Is�2H�kg.~v:�&�2�i�K������� �+h��r!�����A�T�"�^�>pl�~��3��m��h����8H�[D��K'�S��搇JaG��x��Q^��p�i����Do��
e��2�~ƻ�O3��U�t(|�a`�g��V���7�x�L�'xy]x��A�e�MR,�������c��L���9�ؑ==�Yך�7Q��N�`�f�S�$�>�����Xx�`���I�s�����������GhK���Q���]˙����rF��Rs�ƱMk~�K���s=�W43vpR��`�6����gp���%�l.�>Ƒ����j�qxX�矚]�v�;><��/O�B�z����3--�˅��Ip��4�4RSȕU�/rg#Ԣ~��-�����A��w�5}������Q�/�bM�����	�}v����dT��i��i��UC�>��R5Pr�mf)3�Yo��w���ۮ�qA-������j*z��Uq�D���׽8Ԣ��=�pvEp16Y��c|3Ah��
b	���pQۂ��K-��Y�J��YR9�4T�[��T��GT�5�s�l�d%cu�쮻N��Om��tΏ����0���>��j��d$@���Y!���Q�N4o��d+踴�:�m�v�$����y7Z��B}~]����D�obpG�:��ye�F*ąt7J�,��x�8�����:@OS�����.U��R�l���,�p;N�QS��h�)n����%ʵ�`�nڊ����d &t��L|������{8�E��D����Ny޵��K9U,@b�5r�����ه2Щ:�Q3ĝ�=��7��?����@p�O�](�������ۊ.)�һ�I�7cKЂ�����������3�>��,���7@uhH ��[��b�o_����.C>?ty"|
p6�"�Uӳ�DL-����>S6[i�"%cu�eY��C9�X��Â�%���,�uӧ���U��KHl�J��$����t��̙�b�ѧ@�w��+�'_�w.G|n����G���=p���]�{���lZO�]Ku�^g��Y+����G������G�C&kz��k}־����|���@pr�Etݲ]��� �H����bä͂���#D<�N���Z�E�"!���D�7�-�uk5���ɚW �u"S��N�y�+���}S]��a;t��g����墣���k����c&��x_�<��X�y����"��a�{��'�l��:T� ��6;<7��N����W쳢��H��'�Z7����;�=�sѲ]ٟ0�Bm��hT\ϊf��|��t���;Ƨ���z�\�K�����-�I���D�9D'�~��ک��U? �B�\3� �t\;��v�R�'�+�;��G�&�6I�E&p(e�Ț�w��iТh��۹o�~�+��R���]i��x�Z.�f�d�N�ֱZ��1�&S�Ԯ$��(Z�F�����DZ@	�G��eI2仺j�o
<�:�J/�X"3;<��R+tA\��!����9Ulf�I<�<�m�[1u	��B�;Kk�/c��p:[D87���3�A%J�ZIV䱺�#6���X��/c���gJHn:��!IA��5��R��f��ӡ�J]�O�pO��Z��;!O�w}��[�$��a��"@�%���� ��8U ��fEj�:�[f������o���G�pO�Q��^���'��H���N��6��G�I-��':A�\��m/���F��T�}F���iB-�G'����'d}I��_ܠ�RP�O Τc;�e9H�����1g��םt<�T.�%�I��(C:� �M�-��r�����e��5��[g����j 1iZ��skj��?>�u�Q�: �9X�$�߽�t���E��\c�u�2�@�W
7]�����K���
��2*�9�gh0H��GH$�&���5ͮ]M1TZۺ����'Ѐ���ZM��H����:���!�A���W�9A	��Jn�8T� ֧m9Qqs�{ڷ��;!�I�?Xk���b�.~�=���� 2�~�/I��D���h=ߵE,4��m���]aa;X��f��Ê�w'��!���/��`5_ލ���oE�˶
RAΐ�h ���&��+�t[�H:�iʛ�������/|�'�Q����
�F�>+��g/3�����g؋��j�<��߅w/�L�Ɇ�o�4&�lJ�x"l��Dھ�0t��ࣁB�
8{�<[�B+���d�g:��T�����n|��RGBT=�ց���E٭`#g��Y���ѷ.���y,�wG���l~�'�s��$0?�h������d8B8?,e��Ύ���7���iw��o����B��՜e�㕛A�e���F�0X'��xC��1 ��퀒�w8��i�~Ȥ��PQ�-�� ���
ksA����E����S��拏�(��>��Lj**P��B�_�|%|�����B��)�Gw�1�o�N}���ϰ�Z��w��!U?#��BƼƃ��?c5WH��3�h-c�ì'c "�47�y;�A�t�ö���Z�#�1��e����nȬ�5H�sykI}�$�s�2�����vÀJ���=3��aד�����*����Vz|���s��t�.���/{�����9V^#>��U�!��q���s�9#���ݠ�����������T9�I}�	��3��(�pe����L����Cs��`fx5���P��Y[�%67����آ��zbiPI��B�;R�E9�Z��!�b������|alSS$��2�
H�VH�� ��13�*�o���;����4cQ���,������v0��QfV�����s"a.MМ���Ob�Ɲ����)���xkvQ�Nvk�NV�8v�GV���`����eb�ш9�46ݹ�!��:�zX��S��c����h��@y0��hO�#R���*��u�O(rO�fo?xXqR%ʙfSC��O��h�0�&�c#{('���I$���������G�0��^���HqI2u����oc�Zݴ���(y���<��W�Ҍv%�~&��jlp�^�}b���-��ߌ�HX�/�lBuq��ܷ¶���J�kF���-�&F�PM'DQ���V�����e�2wz�P�}k	Q���_�Z�]!<�ѓ���;D��{��$D��nv4��l�K�x��U�3Zw\F�����] ���)��5��X�_�����a�����������>D(2���E���t~ذ �b������w�:���跳ȥ��7Ӱ�F(ɫp��jJ�����.Z1"&�<��� o`u ����zgO�.qn:ₐ�V�d,z8�E��w��F	~s���[�\�?PӎTG��1���籏�S'��zǊb\�	w
���Sᖂj����<�������a�k``��{�3�Pv�`^&�������ll�)#*���
���l.&7o�9V2�q�V�P����u�"�f܂B��$)x��|&��r��e/�y�3��$~�ԴQ�%�	)���.N������ux]t=�߸DO�ڧ��䉭,{~O��^�*��{a���f�>�]Ajy���^CD��Af;���2b��z;D���ĝ�h%�lO�}!X�v�CS�Jas����k��5%�,��u��}���N���t1�|E�:�S�����푎H�ӭ��6R�['h��zĉR��GW!��G�Ҝ�]ɢ��Y���w���jk�������o�Y#�H+�C<����Rԭ���0�t�Y�6#����B�_��{1	Y�<��r�A��VzLt[�W�,l�����چ6�ԃ� ���$��=vN}��n�!gjL����UGL���b ��v9,�OD�����;eM�)�	�+DM u!oᮩ�53c%��2�B���e1�7 +1=D^�/�ˡ��6��ЅU��FL��� ���-/�Gc̳�,�w�3��")�0P6��H[۹n�c h@	���K�P	��ٜ+n	� ��_=�Y~}\�×l.�΄(K觬�R��}4�qǧ�t΅�'�rl�9�M^���yy���b��P�2��'�]5l߸�wV��ׁ��1�ޤr�"�/�+<�ǵ��<�RHvu�R����v�n�I`a������o	Ry�چ$'o~�o9����VQ���_m����e@/j�D���3���gė��`I8º#��%]��Po�?8-U���!L{��-dFW�o��s�&��KRL=ϯ�u�`�y�����y-�	��x����(��"�	X�y��x5�m�L������(.�r�I4�^��tc�qx�FQ���УhY�^=��19c�>1r"�niǡ(��<;в����6�� �,�¿�ɇN�ˊ*�*u����a�ɅW�,��w�V��E�%g�(*2������1��4�
���(3S�8�҇}�tԄw���M!���4��X|�Ӈ�VsI�I�؝�6��*��p�|��oWWR !�����[͢��#9\��n�¼cc��Y36�ِ]��dqJ=�>��'���	2)���� o#a:$��r��R�͛
�CFrڦ~^��yɹ�&=V|؆5J��"�H�L�H7��{��Cy4!u�:D��|��a)E�A�[=�.xq��~�W��hAE�k2���R��P٘��
���o�u�����}s=���Q����n-ᚧ���n�ؾ��_����`K�!c��Qz s"���	�0�a�� �##���Q�/��������
�ۈ�5� 巄�!�?,g�si�&�.QW������ ���&L>lT�j>8[	g�W���8H�W[�x$�G�P��t�h�����cI��X�=H�v�Nv���w�nL�	-Ԣ�U	�;}�����B�����=4�B�Ĵn�V��n�?ҳ!acú���H�fg��;k.����4;C���� ���Т���|��/�����
���ӟ�Ғ������6�ɵdx�W�.�շ5?R����s���r�+��@To%9؆�3���ԩﱤp䨊��Ό`�[�b9̟XD\"���؈���
J\�U�ґ"'�1��PG��~��2����>M* ��k7�aaΥ�r���k���5���d o�us�C���fK�vQ?랚�	^\�k��P8�����uS����TT\����tVG�@iӪ<wK���5�͚��+�3G�.�?��T�����A���J"D}�5&��4��HE1'n�P4�UkP{tdw$�>%g����n����5�C�醴T������G��P�,���5�AN�SyO�+ҷ
�9�?�Ğ^ٟA�/�W��߂�2����$����oċ8��j�¢�,��p>�<�e훖���=�^k��5i�su	$m��4;9����RYQqp&C�j@��1�xa��O8�1 $�y���wp��(���!�ݷG�`�5�4�>;���k21��>]z�ȭ[}��],x+Y9PSc���iL�9At8�7ť��1g(�o�:�w�w�#�7��>W_��A�?�Uw����΋��ȥA�>�(���e�-�A�;T0������EuWpP?2)K�i�&s�i��������V��D���9+,�0����������/W_������1I#�~�e����k=q�k0+�č�n��1��!ȯ��蹡�����K�ؑ}�N�������2�B��|�=,�a�x¨W"��6(*>���{u�*D#�)�� �z-@;���g�U�_�d?���l�dq��Y�Ո#pӈs�\7Yz
��pⶆ��KQ�t�����8Xa���l��l��=hVL��(���n�I�W�˶��xڞ����M�IQ�����^��{���tߨ<�h���T7�숞}�[����0R0���M��!m�<j]�b�(ܩ�_�s���զx��'��|���#��Y�TY�#��o� \=�Q��MV��!�(,,_U;
�{gƃ���z�����u�r�?*z���x�+�&pu���$nj�X���O��*���텏�U�&��K��~���P���{Wd���W���M�bRzj�pnD���q=b�Gw1@��trz��c S��I̥P˜�_`G�=��=U/'i��z�43�Za��:<�e�ج8J����"��w����%���8�0�Zu*o���,/��>��`��[�Wj�vy:����e��u踿���H��xX�Y{�	�K5l,�_����~��s\81��Ԛ�q?�p�[�-٬��v��b2۾)v|?��;?��k_�yG��HQ��Wnw[�ws�
1�(��ٝ��v
�P�$��&��I}g��F����x/X)v�w��$�u�N>�j���<�9d�߂A��"����s��Mm%>Bf�vV~�9�z�����Ya��j'W�Жs�DI�C�9J��_����GT͆�"�V���g������,є�[��re��-��;Jy +ݲT�C��y�Ѐ�ߠ&C���
��)�$xD�i%ty?��ĳ=���%p�j���|��x���k��#�Cf��O�6`��
�G����7�W��ٞ�D�� ��6�z�[[�e5R��A��d�K��U�/�b�W�S�S�H��v�d\�N�ikO[콚�\'{T��~�"��u%��z�鯩HQ�#o4n�ǫ���Qy�W�����kc�.
�N��h�UÁ=�n�� � }���Y��
4
�����A02G��(e��Du�=q�g����o�%%�:�3HGo��_)��.�X!-O�$��E�B,ë<m�u_��)p/M�45~�-�ϡ���.<���lqt������� ��S0~�6��l��
=">�I9�'x&�n��y�x(�I�rD��^�ڲ��p%'��$���D�n�m=�Oo�T�&�6�((GO����H{�/Q�P�v��/!���8J�yO#�&��y���J�xH���^�aT	WK���T�C�Bܜ��iì��9�@.�8�ֳV%�y�ʶ���R*��I��](PK����
�L�+��~2͙֒~�I��7��	����c{�L�R�=0�y(~o7��(����1?�ik0�K$V�����R��Ħ�-���r��>���?��Qx�v[�_��	P~���n8�(�@�6�}���0C�{��I���T8��0 ���V��i�G��˙�Ҵ�"P�#��?Xe�[�2}�Q�Sp����HuB�xU�U���ѩ\��'�6��>��P��є^NR"R���.,$i/��GQ�BN�Q�{�yC�?���j�5�dvT���L��1=�[�^�p�;ZW����i������K֕��}J)x���7�?M�w�&�����@Z~���1N#�O��9n�;�ߣ������������==��r�[ �Z�d�
�/�ա�åa��Hj`Aqs_�:n�ILm�c�5�s�h��AQ�Ejx������f�)�3�"��W[䎏�A��[7x��+���M[�cUdy��^-@l/��׭��=|�<c`v;f���wkC�nΞ0����lD6;,؈Z&l��g����n��Y!%��Q�Krx���EW5��������~��Oh��f١ɖR�^9����W��guڔ����n�ฃ2��c>��I�M[���A-2�SG
�'2��q}��v�Ӈa�ߔh0�:�f�eȜ���4�����d�+l��K�}�H�+*�g/����)���>�ͩ.�9��˵<����EzT��M��׹��D��d
%8�r�tV�ZK*��`<x(g>�(�N���|r�Ӷ���Y̌�(Sq�ׅ��8�w���lAFC�<"�k{�J��ҧMB���Y�S�|��O�hAA�%=�Vp�l<RYo���\���6[˾��H�v��H~� ��kȎC�S� �γ=$o@��{�1��ȘC�(����B.R�������v@Dͻ�z�d?�M%l)�®����B9_�y(�\�yW��IոWx\���UD�D�b�=G��k�a��4C~�|�U���k���"�P)�x�V�\C>`�螅颓�']@�{���_~5_�m�Q�J�y��t��Y�q�c~�^�"���hQ��J� ��oA�e��jTȢ��ЯU@��A][�]�y�wh�\�V�#Ư�/vZ��DK�P������7���0��rpj��I����]/?��&�[�nM��<m���cu�:2*��H�up�,4,l�1݇�g�aZ�g���Tŗ��ɇ#���g���[�Fۺ1<˱Z��$�!���5��k���A�w�O���̎�SyE)���R�đ�e���WR���4�[3Ά�To�.h�q�@��+��֞�)�l�V�r��bp�aP�V�A���
�J8�P�~�%~�b S%�?�t�*��o�b+�q��..<Q.���[�u���X�Oܞߎ=t�ؓ����#B+�t;]�;���O�.��|�P�jE�{Ӷ��_f2�4�X�I��c�<!�RyH�gI<e����p)�Hu�j 	��_o�Ա3��	������ah��T�L���ዅK�	���t{��
gs�6D�,/�WŅ�ݸ�e5� �����?�^]BA�,��9՗�Gt=�����#��^Rp�دp-w�k�UV�.�NY:����'a�����"�J��=S��Cdۄ��^���Eۊ�߱������X��ẋke�˝g�'p4��$vu�V{�q�r��;�a��5u{�E������Q��	b$!�`��(��5��e�#����rް��d�dL��F)k'�n�@3�HM����q�(r_��i�~l�������z�E�[�dk\~6R�Kl|���'?{�_y:I2�q]j�&�>wGb_F�U�1f)�Jc�>9�@�v��2:d�n�z�	��?�;�k��������T���?�RbC�M;�9VJ^��g��J��_N��z�H����q�NƋ���1��p��SQ�9�H*tTI'[����t�QTN��Q�V0�w�0��$���?�;��C\�<Mqg���-����?) ������P�ɭ�1[wrX-�t�1lӣJ�!J�KE4�UE��5�r��"-���4Q4��SHX���@},l�[���}������競�X�0�y�y)I^NH���|�;��[|W���� 9%��&ܨ�x�3����߰�'5ǋ*J\.���56�=��ңsQ����\RV��1u�9o�")!zCS�j+O�bX�83��᎛|5U�=-V�_տ�9�Csl?�=l�����(fb���f��#J��е�4���L���N�9����_�X�]�,�IW| ��iR�g�ɀӜ@���^G�/�Y���W��\=�c��a� �_�����_�&�z�q �V�!�����Q���يp+�pԥ�Ɋ�?�Vjc�����-?����x�w�5�8J�r~'�K���g��ԃ㐃y�����X�Nw�dvyMʳ�iػV~T���.~ .�&�/:H�<H��	�DQ/%�G����"=RC���ٞ���,b�`�3�ڱ;U$l�� ����Iީ�A��	xwc�����:����0��6w`���eV�s���T;�	�k0����k�8�����A�\��}.j��o*|�N���A�#b�svq�%S�#��K8i�y�J
YyXs �5Ya�E�5M-�v뜂��^gn�=(DTs����:s��Ѕw)[���(/J�ҏ��1/WF�m����v#{�ߜK�2��7���Bw���St(��z;UG^4���t>k1<)O�d2�EU!�)n���F?p�+~f�bJ>.p��;��dCUxr�����Q�@�"`qVWrx�;�¢:��2�hqy�Ü[��+*��t1ɣ����6gR��H�q �@s�U� �����C���2��T�4i�_����;Բ��|%�s�>�R/�Vr0w�=��[��Z����P�0'�\߰��.�6[�B��֠O��U&/��Y!�16�~Va���\���	Q���n^>�ŕ�!��b�PR�kNO�J܉0֓啜��0���ycX�]H�#�lK���;��Iɏ�-�[�����S�i���N��r�oĩՐ�����GQק��^��`V�`^��k1h%���M�_}�d�0�1����K�vS'Ċ�ń�n���~����ʍ�1n"d&"�E��RBE2���?8����'#	�ì0v'\[�_Gf/�����硟�@AMw��^��n�aU�J��%-��5��������Cz=pD��M��芕�����NJ�x��8��<*�Ԑ�)��+�F��
�x�'���;L���i���\Jr//k������Dt�ո��Na��Q9�����<��X�x<z$NA�~a���H��R�ͭA���͐�da�}\��O�Rh��+fL/]��������/W�_�Q���V�Ⱦ�+1ݼ����5�rv���@;�Q�&TX�jQ�}
-��B�{����ˈ;١��ܟ�݋"B\���>�I }� �| 1��Qk^����6��~�@��%m��e!�,]eXM�Lwww�Ń ����	�܃ww[��.�;7y�;���sNUͩn0E����M�E�ͷ�{b�z�/�P�j�UD�4Df��\���O<~ǜ�(��6Z|kAb� gZ{,��:���Q.��ܐ���QM���&|5��ĹcI~��Z��oڡ���8�,��1溾R�	�JM�z?[ħT},��e��(9�*�E��\��>�K�u�(no�gyd�W�1}�\��g!3���	��\�	^o�o�k$|���NLߩ��أ���xI�����ԕjڙp���w#�'�ބ�9�'������&�_W=�D��_ޞ���EY�v1�Ң�l��)�I>WU?�O�#��D�W����R�����C� (�پYi����_����
}�ѱM�K6����H��.A$��s���U����2��;�~l"Ϧ�gz�g�y.��۴���VD��������*:'�@$v+�*R.����x�5~r��sNq�C-r�|�Cr��*v	��V�w��I�!b2-�G�`W�)�T�s���ˈ�A�^�naz~ز�G�s��7����O.J�K������,1����!���j�!�&s�����ڇ��K��I��]_wɎ�J�����>N
�Tl|&�%�����Sa����=;�L�&E��J��&:J��T7��v�J*_�ܔ���f��$|�~��1�(_��Qҏ��9Q�tX7��fWC���?�Q��0a�y�{g��QD"1SęS���NX�co���`[��,�x�78e�r��k
Z�z��Vٮ'1֌�do6�lL�И��+=U�&K��S6�JlЦ?H?=��+�������"��y��br�I��G�¢�����*����M��i�����p,blE᪏�fY����ևQ��N�0e�:��!ʈ�hA������fy��CaD����h�b6�E��(��j����
�Ua޵k��5 )VYfl��F3p۾b�̓~Ia[-�Q�=�r;73�aM3s�W�g+����ƪ�~�_�:3��ݢ�f��[X�C'��I���k�"/YC�YVO��q?(a��J�W$�Z@^�g��spU:	6,�ZI�S�q������v�����=M6�>\�+��?@%�&� &�.�F�l"�+�͖�+~��}V��
@��d�I���%G�i����ϔ��4��0���eI��}h%��f�9������^�bHY\ZX��s� I�پ�������0uA�6��H�Ƚ�wU��O�o��Y��¯P74^�\���ES��S�g%���LﰍP��mگ�E�]:Z��(/yGA�B�㼿�5H"�N�R�U�����іo�y__3j0�[\��5+����$��K��2�R,J>!+���-��Z��(P3N���N>Sⱙ���tL�.l��GE�/��[�qtk��nV�̴݆��9���CY-���3z|ʄ"ț+���a���(�p۠��.�b)i�����Uo�?�Ze�*��^@����@��v�@pz%�M����2r?5sc)#�<�� k�n��T��=�����g�)ʓT^Y�|��~ڸ�O��h�K�T�i�r����NFm���4[���$X;n�l�e���V�R����!�F��
�]uIU/�pt��x��0�= w������/��
3~����'���?g��a��?V;�Vy5��BgJ_H����ܢ#�z�v�mk����'G�ě�[�z*L�^��)5��A��Y����me(�Mt��S�$�7���.�T,Dl�����JY�%<݆�5"�Vn�&���p����h/��Xz0�W���M�!�0����l�{�_��	�B����]�~j�5���Y��<vl's�+���#ZLp���wr�*��!����uy�y�!�6�1��4��d�c��'r4�eE�
��eA^��2��1�HK��r�Sy��}�u��؟���M� ͻ8�x�Mc4w ���,\��Ĩ?A_�(G��,x�B���d4����}1� ;���~)���){�[EcbȾ�h�f0^7T��G�mR5�@Q��m�^��@�o�o���~�H�I�z��m��>�&�󢠪����q	���*��B�E��Y��~P�"�C��k�UWF��a؜m�|�i�AX���Y���\G6��R�-���� o%S��b���\s7���O^
���˻>a���(]�
ju�Q?�vos���1ʴ�˭<��K��;��m���L-V��66f'�׍��B!Γؗ|���w q�°�%/���#���<�@�\�n�����~~[l���4���@U���:z']�����a�W)U큦ĥ�m�G���F#��^&K,�fbLa�;�˥�T�cO���i�T��b�a)-xjG7����o;��*�_������c��~����������~�߈'��>�;��}.H����m7ҩ,TA�J���ݴ�x�W�d��ލ;��=X��h��u�F�@��?.t/@e�j�6�bO��Bi�"O���q�wN�>��<B�������aC�dr���ql9p�B����H�">�? �2�
���ڮ���)p���b�W.�e�ł�w�f��Y
�\h���̬qF�4,�#�|�����&1F�f ,n�y���8��9\���s:А:�"g^Q.�;���J=}Xws��m����}�]}�ذ*� G�f�$d���e0̿�gP���d4��f�r8��5��'u������U�e;҃����Ӛ�A,�Eu)F[��4�H���TL8+�Q���?���爝_�(��I<6�{>��N`V {ܭir�o,wt�}�sq=�N��
�^�ǲ��//�{�_�^�Y��h��ҋ0��)4���. ��t���:!�&���}��/�xg�a'�on��Z%��4��|�
��љ�֌����+�ɰw�f����so�'��r�t�5*ꇪ�@֊�d�%�]��-z�m��=@���*+�D8[{g����nب�s�Ƣ!ʄ��ز>�軇a��tC1H�x3?����U���}Ⱦ+](��[)S[����:�k��$��2��fk ��b5�a����j1��N� [(�"?x�G�S\���<sYut��).M�f��~ǹ�\n}�ɸGk-�nICLYO{"i~f<Ja:˪-RF%���@�k�	j�7�07��67`�K!�b!� @8��$pG�;�������s�=ʋ?�A�K]\j"�
��9_�>������!��v�ȋ�m>�̚��(�?X$��2\��.�eR@8�{�(i�UW��O�F��ȉ4Ņ+��Q$D����O�Z2Ƌ̇$2o)��]��I.M��x��x��A>[�o�d�C�����U
��?-�bA�UZ3T�Д��6���g�%�6(���D�F���L��G��dтk��.@�VM�W�f#��$&����`  $�I�l�&ړE���rr��wV�t��:6�r�n����^M	g��p}����7h�;�4�Q��.l�wϣ����Q�r��^&J3A��"��
�\�G�~L�a���#�])q����6g�/2��KCtB��ts�x�4�}���
�Ң���{���}��β�����y
�<�OU�K�j_�HX�w�D��Pǥۨ�j�:;l��S���Ww�G���7fЩO�.=�8I���x�Wy��&���x� �v�w�����F�bMD�iii�KTC�x�;n�a2�@���v1NL*��[d�V㡣��<}��t�,M�UFC�-糀$��TnT�$δ��Gd�(OK��(�A�q�N��d����a+��5��4Q��6�S�!-�U����(��y�P����֤vɈ!ٹ��Y��h�h��-�n��tp��c���=]c��e[�7�l���l�$�t
Y�y�,����`R�y2#,�^ћ�z�s�����_�R��b��\N���=A*s'��-*?M(i�ಢ��ֶg B�AN�񨄵۵����;`C[`�a���n=8Jw{4��LAӑ�����/۝��`/y�[��J�Ԉ�T�@n��24��nxw����kѠZK��E
���<�g�e0lw� *��L������Ϳ�j��-��p�u]�	%��pk�j��_�wۦf���%�BS��&���եs�4���n�h�\&��-�^��,�:B��"��I{���m��0<?��3V�s%�n��f�6���'�yk"��0�o_��{�&y�:Vj�~5����!?��`��N.�eG�b�2���Z�����`	w�r(�yq��~�<q��{����X4FC>�7��k��+O�'�ί��a��ڕ��t��
��T���ć�!��pj��+�NϻS:����^i�9�~c��'�F���!�a�4ј
��X�����E��я�g�e�/��2��u^ގ�xCN>U��a`|{�x�}��`�IP5#�bm��ˑ;�惡�H8}ĔW��)����;K�o�ԣZ��C�CW�Kе���#Yb��C��E�g��:'c�i�I����_ i�in.^�b.^O�P>����ҕv����T���I���B� ��,��Bi$��z� ّ�U����ؐ�z�I�r���s���삚6�y!����UvԊ!�C��\�?g�)�ш^b��D	K�Y3����o
��������b�0��.˧�"�%Rr����zE+<8n���1��'�����}jUi� �I��@_SmS�=�W����\ݮ���s?m��a�}��li��ѧ�I��3veq|�Vl,. ���1t��G��Z{���P6�Gў�-��h�ny�@��b����`~�O�u��x|pf�y��?�QR��!�����|������e5�]�[���T��������f�oU�+F���mY�Rab�K�޹���{!�E
9��"Y,J%V�1_C�E\@Z5'`[��r,�z���8o� h��H�5�t������_���� 	uJA�]����~�����c�49��/T7/E��f:��b����ؼ�K���ӪF��87�V ��~��IHq�YJ�-�\i���
�D���t�ñ�g���X�l�&�@������$ɒ5��Y��� �J�P�b�<��IT�_�dI�J[��y;-��}W@b/JA?6�[�Z�ɭz&?B�h���G����ԥȱ�pu�V=A��W��ᑣ����9��bMsQ��C�(� �
����6� eK�u�j�od��O/�df'�ƅ?�8������-��]i��@�X�s�47|�*�gجqv��Z�S��_:����W8����g?�RT(�F/j��h�e��TP���S�����q�[PO�eݣ[���ei��l>���|\�އ2L�N����'6�EO�?!��tuFK;�h�R~����U��O���~iC���EXk�+��BHC����.��	��n�&��i��GR�q~9|���H�2H����u2h��Dqc������U �¾�E��񛯑�d"["�^L�����CkxJ�r�����'ĒK��G���!��pF�g��;��̣���y9>ƚ9��bnA��;�����ƕ����R�.c�f��Mt�h�H0L�P�,ԓ,��"�S#-���u� ���������k�����[��VLQ-}D����ȁ��,�
z���[�É�{7y��)FGH�5��jF��gAyQ6i��Mm�5� ȹĞ
��s�KӾ?t"��k�Ē�_��\o���5��l��,}/E�?
��+=�04*O�98t��'5��gD^�h�򽈅3N�|Z��LZǧI��&���ߊ)Q�rC����nݴv���K�gǼ���i�=�ʕ��'1�^:�?]v�}�B��X:�)�>�g1��"��F��kaV�հo�|�K�%8�kܵ)9�:m}�x#fF2&��Ye��7�B���+4S���g:�+/׊�j㚏��I]�R�GEp�R{G9]\^�@��nQ�c�������[`*�4	�캷���7���n,�
fb�Q�����C�����q�,��?ʥ:^<݆J�`��K�HN���`�\���O���0z�V��(�|j�Ґ��YF{��� Da�h:�5��,S�"LKB\��v��I0E@��e�D�D������G"�C������f1W!#��H[�;눆2������&�������d{@L\�UZ���ӼS((��H��J�ы�w�Y]U��'�M�_�BV}���E���,rWL�d���Dw5\HqUW�}����h�����\�u���'[Wi�Q��+L�'�m9o�LŚ��^X1�[2����,��t�?�M=l5^R¹���اd0#�l��4�M}���}�l�Y��(qrc����5�B�Lݶ��,E>�1����$m����i]9Zp����w��xI�%�I)R˯�p����\����ۊ������XX��F1g�>B-[�Ӕ8�yv�  d������	�&���.Q ݩxv9�^��^���U�,�W\��`�V����@��!�G޳�nk�s�y���;R��V�iݯ+���R�pP��kw�6hx�\��������ȗ���kv�������I�SojB���!w*	�M�C����8��#������I����\�`�78I�*�=2�"eA3����/x ��(���*��f[�v���,Z1�)d��9k����h����/TD�K��sL�G���0�w� �hn�s�޷k~6{l#�Cv�e`�K5�?�2��7S� Z�^�y������a��ײo:e� ��l�U����s&��aƋH��n���r�j�v/R'�����;�F&� Wd=�L>gl�?
�9����/!; tyJZ� W��\f�+���a��˟�$5=���ZƤg��M��_D[�r>6ct:7��~�
I��۩�ԗD��
;�a�������b�J�����F4s��6��4����U�sz9�t���>h_��~�ۭA����qI4�"u��b�s����<���gɍ�ߵF'Kޅ�0�xM�!p��cĀ�I�[�ܛ�H�KS���3�2���*�S���31��o}-M��}�6����Wm��x��R��>��qB,�$	�a��wP*+�gtP��/�.��0�1��JB��l�I�:ICm�HU�m�z��B�3�+u-�)������iN�����Q�i��|T���p��n txZ�.�~�������(܍<�bcЏ�%�s�x:�����-�,�	\�C���R�{�8�;5����bo+��+��~{�z爾4w�8P������dF�#�gA4��cB���Q�g����hBHB�E�F�S�gC��;2��_�'�Z�߄\�V/XV3t /�UXD�l�`Q�e�쿣"�չ� �m��,�*s׬p�4X;Q*�M��T��#".4W���V̿c�p>��]�Dsm��*s'r/��Ѷ��+��T�-���ȓdR��i�D���'�O!�d*ҿ$9��i�B�z<�(n�Ũ���cLwv����1���>n�A<8(��#ui�#�2�s�]��x��0�G+\��wO�9��Hx�T�����p�� ;���	ĭ,����PK&���)�1V�ĭ��K� `M�N7u�z����tȦ���/RU]T�ٌ����(e���n� �<����?n����x3"�w�D��k]��#7̓�[AA�+Bە99�������c%8�SN�TC׼����]���}�f��� ����#F�c�bY~١`�KH�(YʉҮ�_��V�tс<��Q|'^������/��H��a�[;5.Z�X�f�{
|�E�%D`������G3��m(�a��C�����8������-#>ZO���δ�'�����Bеو�5!pmK]J��Oy-��Sb�+l���أ�/$Uq55h Kmw�Hu�%�Ë6��t��rSw�5�hq	�x�&0��KXy�h�L��'[f@#��j�`E����E�+lӬ�B�AW��i�qӕ�{�{��T�sU6�F�9�,�lYA_�2e�!?�o"�����<C}��Z��O<��8������c���$��r�>-OU$G��K�M�5Y���67�B�!���]C�|+&;�?��������L�;�*�%�yoV_ �>pa���bz�Fn���pU��:i��X|�3�$�%��V���f#��
�B� 64g�NV���i�?���,?���;7��ٷ)��<d��M�e�mw,��宧%X����v���mX�ʢ2B�V�5�����>���@z�≜.pM/��C�iMq���p�أ:E�)��ϔۇj�y���W��}@Ź���y
�6�C�iMW���y�_�9�'�Sv&'I�<�)�^�3�[�tQ2o�z8Mܣ��pߠS���Pke'�K@{;_��[��K��<Cf��-x�'W[-������H0{[���D��FϨݞζ�)Cd¹n�H���JϽ��Sy������E�K�?�ꬺ��:�E#AФǋ����(H$s���
����P�QE�~��D���
�<��ٔņ�pDs2e�R`N	���+��r\���ͺ"����ҷl5�	�������KtY,ǲ7#S�t�1�JSŦ_��L��6`Tz��R�Ա��쏑3��j̑�2�M��s��}g�V>�?�P��"e�NI��YH]��b���.�zt�,��h.E��f�i*�.o� ǈ�p҉Z$Ҏ�D4z�*��X����S�t��Wso����	����I�9�I��wTN��v��W��p����ѩ�<��[G=�g����#6���
2��| �'�D�?�>M�/�#=C&r'���T��/V+T��˜��R
�,ڟZ��/%���Ah]]R����r��])-��Z���X�*z�0'��ۜBe�C���
�,���e�q��}��?��ʲ([Z���I�q� �)�6��l��V��Lh*���)$�,Mh�a���_��"�t�6��a9�����&��-vxM:F�w*�<������yA�7���	A[�<f���n?ɴ�i��7Sd�x&���ԥ#-���cF�9a����e�|
2+Pu��˷tPڴRѪ�Ԉ{�,�+��pE2k��~?�{-�T �7�#J�2�U��o[��y�������g}��r���>-l6����0
����m*1�K��Ea��%#Է�z�����P����r���>.dk����HZ��%GY�����1�FU��E3����ނ!���Z��e��1M��z�Ej�>�+�ؕ$CyRT��o^�8��wl^PD�(co��F&�Ne@����U���S^����4L�'3�x^��#�!�N<�Çnx�0Y���-%JμQ�����{=*�0���g�?���ط:�Z0&�TS��8W��_9���k[��e9�ߒ�E��B��h �%���7�˹#���N�4��ˡR��):1��xy�	��E����ל�ER[�1$M�������E\������!e@I$��������c�Y��?E��6L�3_���i���G#�ok7l��`ܼ�X<�g�X�"^4nD���qw����K�\��n|��5�;g��,G��)���:�I���MhE�PS�%o�A�{�]�@�ۘҗ�կ�IiI+䈉��6�̲��M\�-���A�S�K\a�<�A�|9D���#��-���@�m@�O��bݞk��u�t� �����WQ��0�ngc�Y}�ߞol�gB�6}즅�:$�j�cww-�0D��NE$b+����nTma���'�9�6�˄����sX�z&��&�\�>ak �O����\�/���0�ݠ��wa��ںJ���k�pY�#�c��B��\�7>�g��0�j;�;ݣRl�F �`r�$�1�.���%9���7[}��.Y�K}(�Y��/7�yZ����Ϳ5�Oz$KLL����G�[$V)��?��O):6���{^�<��q�����L:�`��'�Xb�nz��
�[����Ѱ~qy���v%2�R�,�,��lG���{��95��f��4���k#�&p-�[���B%h"����%P~���*�o�7,��hh,�V���Ib�,$G {�G���·�����Q_?�O������lթ��|-��:q���:� K��G��c$��&��.�'$�'[<%Ζ�lQ�"9��R���/OtW��Pg��I�@���^I��Ѵ�h�~%֗;�Ŵ���A�� �qj��^�� ���q���@{yA�|+%�6��(a|���
��S�nM�ֵ���Ҁ��_@��HY�.���A�*6��j'����ʾ��|�&K$�����P���݆��!�k}y���~kyVO�M1����a{��k v�+��X��4����Z����	=,Ư0��)��������kp=��Yix/E�maH��;ռ�A�����:^m��������j�w�w�<)�c�ː���h!yT�������hj"��s����C�C����������at_�M�
��h�'ov�#B�R�J�l�]�������(_8�e�� N�h)��~*�q��+��/rgU���5�ɠ�'�%�F�Q!��w�"���?�'\b#���ԇ�pFˑ�k��.u�p�<���d�Z�ov�*���ڡk�S�".�͐��<_��.�IV�,3��Y�p����h��о�t��}��6��}�j��Ӹ��ʗ,I��s�(���R�$
������y4�'�m��w�6F��Ho��+�ޡ�9V��lh���l^�I9���ъP����������8+�50z'y���� }*��Եf�C|�Np2�W�<�[H�͌�C�ښ����Sg��!��	ҫex�g�iF�N�
˚yUL���6�0�{�-��I܊&���su��G�����|�2x���w	����:2����u貍8K�y��Zl����<����K�[)NS�R�&�kݡ���N��Λh]O�����e=�u�` ��k*�T��!�8���VU�ky�qI��t4�k��N�u��|����eq ��7����q�����D��e�����5
;��^��`?#$H�Y��`�'�$�E�q�-����\Mkv߂����Ht`���� ���f<1_�\fN��<@#0�	�v���G�pKg���AϬ�B�c����I��H��o� �Ld������i��Nҷ`*GsB���#�~<��MM��:��Z=̯��/�{t	у�����b��q#+����H鋿��m�qn8�N YS�.�u�eY���tC�}���G�������G+B�:i��碚J�-#3ul�R:wWF��[<����0��t�E�(���Z� p�r+�ݲް��G��Tdu�N��nh��{��L������
�0Y@0*/���wu�\TT����p�9gL�HY��#7w8|	��S���2�~S=\�t~�g���,��
@"@�FΝE4���f�*F+ײҒ�Ǜy�m�}��]� �-��Xu.?0��؍�9�a��L���������\1�����<Y�7��
�G_!���C>͹��$����D��h�h�+	�JS���g��c���Jɘ;f����=��B�Gfk�N� .��+!6��~�ܿ�I-c5�M�J�WE�b�0��m�KfC b"��'�k�Y�$��aC�N� DDly��n	8I!�K�V2q�(ENUts�cd@�ܛ��T2�[0_��a��œe�!��s�չ�s��2��?�M"J���,+a�q��Z��x9�!ڰw������\ ;���š��p
8�/�s�7�Y����p=r�63���N���#Oy���z͚��#I'(^v�r���B(�ZH8B3��m�F+�N����J���ɀsPbb9q�.������>
��s9�Y���~ayx��Hx�`�ah�;҈�����W@�2�%�h:�u�p9M�V�{��u�{���K:;;��x����xZ_|&;�عp�B�ZK���5���l2���[w4�Ƅfƙ}�����1j7?p�n�^���.z��T�Oދ;�=v�u>X$l�J��_4��@,�9ˇ�f��>
/	���i�0�S螉O���kn}b�N�
gTyq>�z�;��v�p'h4�1���TF������.Ui.M��E�8��#����l�[7��Aς���̀�LD!���ϯ24Å*��i�iUV���ʮ�QK|�/D?҂�-93ٛ�[���k�0���U:�z+.o�����'���S�rB.(��Q���e���$B�@�*{cs�V�μ�m��g.�J�����<�SȭG��'�.�����R�3Y�
��&��[w/�SB�"9���q�R��a��@"i[��q���zP��o_a�+B�o���hV>�+Kp��p'����GR�1�ow��c�9�A�H��@�.������4�\�p�Br��n�`��"�5��-����Q���Jo����e~"7���1}S�Ja#�)�Ry����2O��aPW�]8��ləЧ������5����8������D�}|t�'��5�q�*��F;�녭��w����C:�h��̑4>^��[��<9SiJN��Nz��*P����	�Fϭ��H��5LcR��2���qi!��K����*��ǙN���ߛ'(��2�r��8�,��Ƒ�CD��or�5�+8Ȧ�sMQ�1a�ь?A��j�]QY~q�یG��q-T��L�jd�������Y�	�Z��L�c�Y;��ԐS����YM�����F��O.?=�V�/�:��E57G9�j)��^-Rp3�̘:��$C���dZTjK��ݤ'����TK�����4X9���9?�o��v�G�]������W��ЬIp�`��#
k�D����4ѣ��a&��y�\g�M(��l��,��Ա�A3Ѣ�D�GLM3{{��tH��(azӣ����<R	�oF؆v~����� � 0�S�}�Sclq/�(= gl���<5˧���4���@��>\�e�D���58"e32l�Z�I� %���B`n��ƈ���wk��������,���.��|q²=���OE�ͮlh������yAc��o�Z���Áf?��,�-8���
Ao'<�e]����n���Q�
���QF�-�j��H�O}�!=�
�"5�%)�&E_�ۛPjr�����g�r9g->-{�G|�_���r����'h�M���>��M;����th��������3]���E���G��Wx�K�#��u�S�� �m ]�#���zsT����^���!οK���k�O0��!�:k��EޑI���ɻH1d�
ys�(�x��O�B� ܚ��-/Ȥ�=��=$B���yd��ϗ��zT�#�M$�H]�p�� ����S����Z�;E�����g���[�2��!}\�刹#��"p������{�ypi�\Q��<Vc���TW!�ljψ������(���x>E��}��ټFAg9<j)m�u#����y�� ��zP����4�U��ٙ�")b����w+�S_�\LTe��"b��S���,sB�q����f�yl������xݯ�L���`��������>�L��4kHiC���O�����<)Np��?i@-��|�����bMe���r�sĬ����T�\8�|�����t-u�9fG�~O*�"7B��M��U1�2l�2|�#����鲦��j��bL���Q�6�C��e��'��/�|�í����CM��E�1��\`��	GǮ!pL%�3W�i tA�O[������4�H���"�����%<��J�&2�w����hP�[7�ͯn�R�G��d�~#H�V�?����O��{�p����H8�߰�;/��(��#�9�K=�;�K`����8q!b9��{5����`���{�"�O�A.s����U���{�>{ۓ��=����R�.���O��5��R��/ �'/T6�U��Pr���|.�)4����{��?w��h��o*g"Q��H�ji�!�����2�W���:m���`��3$��à[�Cs��(\��f?ᴞ���EX8��%*��7��M���}}��b����"����٭�i�S�h�M���p����S�ᆗ(�V�̌f^�jl��=Bj���Oo�K-�G�f��i��#-o���I�����oZ���9hPF�,�����A����c��<
�y�J�Ύ�\���׆��3��F�m�[�����-�X�~�	*�����(�N����luߐ��j�(�Z��b�%%ڏ��E��}��&W�l����p.W�K䧞,�A���P|�9��&�u"6Kj�0W]yz�Vˏ��W�u�Ɠ�*wz����D�Q�ki����Y|&�ae�OLGt8��y���r�i�%�<G5���W"��k1^d����w�o�V��n�&!]�|S��]�x:�2��t2t�(p ��a1=�J:�x4�X��p2l��p��T������R�V����2���trN�;�V��2��L��� HҼ��ҼH���Aݯ䂐����w����ID󜜟�}�&Sa��~�/�ۇG��7(�^�������qy�<�n������o��4k�#7�����t|WT>|Z���իK���Uc�ėM�ʶ�ylVuT�t�0�H���#�g-�R�!_�4����m�|�*�w��/�ra�]ݤ�:�W��ިP.�Ge�a�`{�ǅ5 ��`8��;P��܋��j_.�~��Z{_,�mS��Nx�u�\Ȭ��DY���{��s�(�Dګ�5^p�\ޯ���d٫	�l�ݸ���W��*�k��P@��}��9rH;��'���NĶ(��1A�%�������#���I�	6�_K�U`"��T�oWh��H���`��1�� �B��0����{x9�r[���ȷ��p��ⲅ��CM� �����2�
NT����8��!��z�qHD|A���4�Ċ�E�l�q��U�{~� ��0���C{m��~vg\���Z���;+�����"}�p|�ן�z�6������ʭf��_�,����P�(���.�k�>��a�_/��uM�p�
n��ߞǣ� -W��Cg%���%zh��'�a��ɇ$1��u/*^%�Z�[�?�UMu�C��+\���5~��%��l��+��o��=�a�"Vu���d�F�{{"���T�zk^��� {�w;�����B.;QI��I��i�W��^n*tF�U�Z��ڍ��-��xi6���T����Rj�N
�9ڏ��ƹ���ֿ����*&�E�-O�]���u%n�#	��^C��_LA]�N_�l�H����eъ�?.@bR��LR��>U���e�E�����yX��A�y��tA�t��Ƙ)���D,��.�5��f�߀�Gm��V��Ud�9ʵ`9�� �X�f�C��P5hY��i�pI0��y��t�5c�*Bl~ҽ�E͘�玧~��w(S�FԈ����r��WZNw�{1���@ �O�>�/?n1��7�F��U��4���!���1^�6ذ;�R�h'��
T�Η`g.He!X���8�\q�#f|s�o�3��M�VW'G��ʌ���r;Ҍ\��;<����f>7�9g�!�O:��Gho�>w"~k�;X�'2aX+_�v�����RG����L�P�T�y��GΌ�a�6(���l�9.���$�瞇"&D��r#.�3z�F�7\Sφ���̲��B�=�6���|l��r4s�j:�Fg��4_�o��KQ%)/;�3{ Y<��V7��j�B�OHԽ��{���ئo�����*sx�Van���Nڈ���:��ϭ���A�f�ϹLR	!e���ڸz��o�������|ݢs�7"�]����^g9�E���+oN��m�$�d���Y�-,h#�U�}n}u���mRo(H����*1O�d��u\T�{���%�nC��ϭ�;��l{���c��j�����jV���41Dy-W��d�P����,
ė� 閁W��3���F��"�JH¦I�޴X�6l����mA/��ô� �)�g���S���ѓx��j��o�"�(��L���IFAs쐀�P�F:�`{N�-�LЦ�َX*�aB�H��@�á=�),q���bΔ��!g��F{���M�T�2��'�H�dLZ���ZR�Z{���q[��4�ͷ7�l]��L~GB���C6��\��; �*���a��}��5�@�Ƥ7'�i֚���"�4��i�٣2��e6��q�b�q��d�z5-L�Ľ�|߿5�uL&z��-p�-M�[[6#O�-�� �]v�mn>�������e�lv�2����t8��u�z���ΙO;s_}n���s��]�ֹ�e�����~��Y������Y^(SdE;�ǣ��?UVrS�V��Ҭ���}t�=5z���k��q�V��j�i���#e���7J���;�|M�ݚ�6�O��<6���or����I���,5M���{a�b���gg}���ݥ���s�#�F��?Vj��z�2�O�jo��||�k��}	�M9��u׬燛R9.��_]P�O�߽��1C7�����w���Ǐ/����K���]��|z�������Z��]�k\�Nd`H�f�\%'[,)o�fuÂ��z����O�Jt�X��`z�����}�7K�+���)Vki.�������kW��N>��5�γnme̷��g����.�]}�.��ғ7NM�w���a��6�5���ϔ�y����P�A�q�������}&��P�1x����sJh PK   �A�XJ���a
    /   images/7b1dbb47-bd0f-4b1a-b2fe-3ae5ceef49a5.png�Vi4
��lQre�1B�4L�%ƒe컫;"���f�d��%"�Uي�0F�^��KC(�Xb(cl#��|������w�s��9�}�=�{����8Y��ȉ   1[K��?@���A�G�7H8� ����w�<���VD�c"p�0 ��A�ݼ~��b���r ��#[�����}�<X���C_�x̣���u�^�������^�#�yI��g���`�i�qOK��#�ǽڛ�zk�Z��^����w�Ww���YØ|�e�sc���Y�����;�V���"�����O��T�h>�P��j�����6I�b�g�Bޠ����{��ѭ1����lG|�9�m.]rp^�h�-����FM"r/�l��ǒ�W�E�F�/ɱX������0#�<�H+��Wp�ʻ��,� wg)�_I{lt񺃨�����S�����Z@�W�XoEw��`ع�F�9o���|�ru0OM�Zf����܌XM$ؐ�� ��������b�#кb���t��޷��h�4�Z�s�$$Iq5(h�#���{C��驼_c�'qk>`wGɂ,��������$u�Q1Nz|�xw~*��o����n���ƗY?��LpF/�\�����;�D�0[A���
Lw[��4�6^pw��@0�����f�������S�wVmYel��Dmv�Z�{�����.�������O�S�g����uB��^���r���`��,۸I���kK��JS���8�咎H*�g+��s��|��;9S�vI����o���K�q�'�E�x�*|YT�%���7-}��(�*�Z�2������R����lv��v�M<&����J=��y'�l�4Py�hV?���2������TS[˿S�U��s��������N%��{k�b�����ޝ�c��磛�p��(l�i1�5��aZ�ܗ��zG�pl�;�~�?�Ĝfm��?&��k:��������s���M�^�g��n�u��ą��g�j�mnt��ǜ����ƫ�]O�W8XE��g��/Dx���-|~��DE�������^7�!C��g1����.g��C�:��v*�X���dV+���<clj
�z5
����B/��i���}742�!�21\+.����u�2�u��Ԟ�����M���Z��l���`���:�frZ��*_�jBkC�`��g?0�L�#�a�=��R�}�SM��!J���y�~Ov�^��W��-Ń�UR\}A�O����+��S6��������O�*9�H���U�x�z��=\�vۙ͝��m,��#tt�h��]���?��!G��d����ce�P���	&��k1�i������kb����Ҍ��G�� 5����$�F�-�V�������u�wǎ5|V�W7ي�n8�Yi��5fP�5��5
ղT���<�e�H��Tʹ�P�������d=�JP"�˵�MW��V�,k��t��G�[�f[���q?��D�Z�ʂ�ъ�`���Ol>*�@b����[�������.=��^���~eHSro��eۯ�w֟�	y���D�0�0���HS���� H��Z��x�t�~��%��*X.�.<�frw7F��
䐐�������z�k=�4i�8v�@
9���~��װ@��_���<5[���NW^�����P'NE�x�Fk���yD����z� 3�������QLn��/���-骂0+	�R`b���@���V~,�;�J>!�=�d	j)���\��I�ICw�#���R�_;�nK���h�\��
Zw�?$����d	kM��[D�B��6����0��IQ��(G��W-����?��a�����!<��Z�ISn)�
^u>BUU;�B�@8��q�H���嫫�he�X�-!}����L���/�ɼ�Rȸϴ�!:3�G�z.�2-�:��3�mD�<�<���S���u���H"O�WT呋酿P�?�!�	ݘ�e?�1�r�1�����mk+�,'+�>�,#���j=+��;x�� �=���:0ש聽�������(��L"ڛl�l�2���BH�ko����@-�����zl ��k�U�er�v37I�	a�Iu�RD6gnHN��;����� �?d���v��Ft+����wz��v�O�ͭ�Ȑ���.H��#�ئ�3V�w;�Ri#�)��,�{�����M�����4|\;<{��}�"m}���eԫ�>�����[�]p��ٙ�<��h����L��PoPfHV���+'�r
�O�p�k4��^!�-�R��Z���ۼ�q��y&�[�'i�
f���\��6R�xkrt�Z6���Gg���*M������·j�t������{����z��t_f�C846UG�u*��>�� �D�kWUL�f��<��1�?��\ȷ��y*וI�R''x	w��B��1�3��n�����	&iZ��h�\��YXX�dP�<Ӡ�Bܰ�A��»�t��z�r7P���G�U>;��u���R)�Ӷ(s%�5Twj��b46�LE@��̦�h��.ya&�5N9��0�YK�^�3ߥ�k��Ϟc�='&H�+��Y����e����PK   �A�X`$} [ /   images/a8bb870d-02b9-45f0-bd60-404fdaa8f6ff.png켉;��?\_ϣzR�'B�OE"b,-�����f�v��Rc�Z�P#$��R�l��3�c�Ⱦ������{����}_׹|���9���������u��;v�Ӿ
7ܱco	�{77��'���������O��X�y���[�;D>��wV;�0�Bk�D�ۡ1V^�;0�YG7g�����Yw/�D���;��І_�����D����,.����? ��?v�@ў=r���>?Ot�8���g�8�Ko��ve{��;��M��g�d��&kܖD<Йpo����k,ѧގH����@5F�G|�X��9�@�j`S.�'��[��ؿ���\�m�݇m�h��Jx۵9w���{�D�c���W��%\[����vn}����ma��������Ƿ}>�cN{��!������	�#�{��.��26��������.��qDSx�v���61H�~���/ڈ���V��|~
t�Kk���!Q츨(��?q6��k>�4�r�K)�TnG� ���*�E�Op�@�]��\�;/˘a�y3D}?��J�������%�����ٌ�<�U�Rb�pT��f�%�\��$S��J�d<�T%6��#AZ���ǻC�zs��0���?Y����z����c�*�9���ޟ(8B}�Uv��K�!���W�DzS�ڿ�¹QFn���\-�-|�&L���X^�M֫�-�d=꼒��t�?�>,�����3�ah�1 Qf��qːY�����)J�	B|U��"����;h�5횇�p���7x��-���"ǵ0�Mø��3j�3��$���6RɟVS ���Y�|䟇e��&m���>.�E�{�.�Hd�Z`����)�E��w��4	����ۦ	h��;���b(��?���3�nԛijiY�7���[�f���ʢ[�M��-o`+��]�S���ḇ)�˨4�`s��ϐ�5��i=ΩX��\��0�żӸ����Kpx��J�e�ztW�J��erC})�� ��s�>��+Ȭ�?'�a_wu޿fg��0�*�{2�as����@ۈ̥/���pK��~p-j��uۖYo*�%H�Ab$rp|�,���6�FX�0��y=�M4n�G�'�s�_�e����>���x�d�k�������f��$�D�����=��_;#�z���c��$w�����O[�&�V�
��?�ݾ��|t���A��U���à�Ϫ^&��A��uص���qX"����
+u&��SJ�V4S8(�}�")�+��i���k�<j�~-�=w����1#��5�E[�ws<7:)e�wmt�U�#g��r�1�jB�{	*C��/Z�X�����V���E�i��Z.���E�pa�L�PS��<���w��C�Q�S޹��G���)!�*u�nˁ7,�o�n���b�:u�J�����f��A��J��'.f����O�-�g��8B��$�PI�7u���;����z�>{V����K|��Zy>A5c�
/g����1�Z)6T��|�/*��,����MD�8֒��9��++�����4�`z�Mک��e}����ќ��CYI���
�Z���ŤTe0-�FY�=8����E�A�]c�uc��^�/#��F�R��kqbi7�jԯW��U1m�/̏��bh�u-m��y���W>-�2�߇	M�H7ڈ�2{N����b%�뜈�M<�S$��r�Ot��e���K2ǯ*�|�í��������'��k�������:��a1�����J�����������&�#�&W�J�(�bUOx�J<v����.��rcqC#ĉ_�E��f|��%�h0L뻸�3a}��a�k��M���<^���~(���`'���"k�	=`��5�����^�o�EjB m��h*��ɡ�{_��'x������R���f�����Zm��f�4i�U^��AT]��!���Q�UZ/E����ÁD�J+��նܰʶL�%H~�;�g��ƢGF�L?�����ť}����ōϦ��?ʱ�c�����d���^������k�i���IL��@�dh27N(��ԿaUJcmm�O��y�w=,0OL�G
��;~|�*��Kc4��M�7n��`�c\�����g���Q���I��Jg|f���v��h���)�՚���mr�)N5ڤ0�e�X}���{Xm��_�ƺ�"��%�#ǚ�a:��$m��ŗa8�$����N�B�z`���|
��q�~���A����ӻ=jić�Q}{s��6[�
o�J�$���j}�~��P�p54�!�3���A���F}�©��S��C���q��9]�OPY�v��r�Y�0�gD�0��gLm*+�`����pS�lp�����I�2�rP	~!�̕ߔE�<F	n�g��a
L�)ݽn��}����B+	e�h�s �u�L�j���n�t<,�M6S������-�2_��+@�p4�Lʾx��^����p�U���q��ҁ�}!��Ya�� �Q� ��ʪ�S�oC������������l��Okx����m����V��S}<A�mH�\���E�ֿ-j0D�:�̼Lڸxh������e�T����Zl�\7�I��n~�b77�N5i?[�SlD���6��$�pJ)�>x�ܰ6�:�v��!�	��J�"fz)QÿbJ��@��N[��niI�jZ�N`!=>��#o-(�W��\�:Β���	�9�qyӒ-t��4��v4p+��a�7/yF�0�#�j�;#�@�_2���q�B�J�Be�p��?4��j��n*�����3_����j���*�~��v���7���m5�i�!�P�V������P7����;~�M~�2=W�q6RkP��*��Z�>r�&Xryk5,�6�qJ�ϖuԎD�z�K��򥹇�+|�XP������HY_�(�X�ԭC�Λ���B0�������c��f�M,;RP����vQ儅�&Z aa���7��F�r�=�Qu;�HN����a���6��2�\��,Iq�5ăj\���n�OPa��)_Ɏ^P?���Iл�CS�� ��n��M��f�F�AJ�Q�jhȢ���1?P(i!2��"Цx
�?��iAH���I�8���5�Y ��a�|�ƽ�O�:�5@;`2,�1.&�M�hh�_��ӿ>� ="	�I�#s��ʝ����������k[���ͮ����ɗ��Y��6(�_+Ps�zuW���k�y���H�'�v�����wN�z�7���5�5����ˬ˰I@�X��&˿G�(�4�0f%��O�#�e1���
G�3�w�8fU�Y�k�g�6��M��m4��'��L����*�G�F��|]��ߘ./�t8�:oYԾ_�`uRRleŋQec|2�=��W0����<&��"��t��I�؍�6>tk�����R�|�U���񧒣a֝�,�^���>_jo�͒��7�� ` :OiI����X�C��|�_>�$��$Ptl R/��л?=�;��g��*��5�
�UN�s(��w�*Ս��ΟU@����+��*G��)���Y�x��%vUލ�X�uS�"X�#'P�O��y�_�r6JB��7x�~b+�)⑰��&�G��[K���ק
f�<�'��N��y.R,�$bΧ��ʬ�o|�:�g`�v�
s�	 �wp��e���r6�Z<�	��34U�_/��2z:rl҉�F�ޗ0IAkv�̯a?�r�b�g@����i�	�j�N�N�?M���_��I�I�KD`Re����3�z���T�����H�@���
���i��G���������z"q���Hni��}�Z�G
�,��)[�=Vi*�W�Oc�*�j.����t.�V���,�t�a��
!7S������䕘�ƨ�5d��uX���y�]Tpd��LgA���`�:xgh Wm��n���g��kȹh������QX��+�I���a�kډg�z0���n-�Xډ��xOh���b��Sa�iz���s}�������l���8X�ZX�}u�<�mpT��监�w\p�Mi>��=R��I�R0��J"U�0,+ng��IT�FG���C��ɭi�i��%���r�9��\���
Ǧ�-<Ş���C}�~����f��|#@v%cBLS�� ��[P�����;� c��=���QS��_|ɓ"��A8��6H��X�^QH��t2�nn��װ��gp�V��Ν�<qh�J� O��FIH�T�<	6�`^-(X����v��V��>�����%�;K��Ò��t7w�DPn��[��ZF�[_�8�������H�\���ݘ��0�`ב x>�[�\�⸓�i���Q@#�C4���7Pk#x����F(	�/r��X�����ɽ���D�j�| ��k �z���c�$������yiܸzE",����h�C�����b�b���D*��.�������[]��\��]ӆӊ�{V�VN��0���5k�$��Ha~��s�ﬗ�ޘϐeW���r� 9}����f��i�vn�:T��in�R[kq��	�1i�|����ˤTN�O��U{u�!{A����w:���l�դ~LҒ��\�� }�!��|\�I��Y���$/�v���ԓ'O�񰱼��kK�Z7�H�W��$���G"�0B���]"Gg�ċ]�.X�;n��6R�{��Q�۬p����G�'��f��6�:�w-��@��>�)iii`m%�^$�\��Bx���I�ŉ�xE�������N����œ�h	�+�>�uJ��D�0�@�}�����]��}ݣ�k����%�A�5j�nq�oY�\��a��Z�8EE�q��u��E͚ C�TV���Y�S�҇'�I�,V$�2[�E:M�my�D&?7T�A#���;�� ����5E&���4����,�;�4�e��̦��
0��,2�v�|���ŕ(6,
��s0�E.�Ҡ�IX_'����9:1U1"[�ն5�;���_��R���u	�F;��uQA��������b��L�'�u�'^�����J�ƀ	se��?E럼!�>���r-�5E�]��h*���!��i�#4�ҟ%������YS����J$�=���'�L�Ȯ���SƏ�
��/.M>}��\��+nll��3�,�=<~�b}u�G�Z.}��0�}" �ɹU]vʹ&�����S�FK�<4���'�]�xXZ`�T��_4��sW�b�VE�2`�b�88{	�T�AS ��Q�����,�g�䔟ck�m��e���P�
m�.��|Gn�Cٰ���TTֈX_��"��'��"JӼ0�a�{25���6�Ȩ�_�2S�k�m4V�[[$c�� �[j�)�m��q���R�,�R��D.�.%{��b"��ݵc�M��_GiJv�j3`}Ȭ�s�T���ӮMz�wԏH�O���7�R�Jt���F"M4k^���b-��5�y�fk)?��Ł
y	��x�{:��V<�r��	�5�>�o�fH�T�H��^6i|{3�,�ɞ�CV����c�T�e�8a�c��d�>��Oi�.�9��=��d�Xt8ȫ	@��a����j��H����z�.`������!�Ҙ}��U�E�1�zfY$3��Ėё�Ƀq���#�'��@��I$��d�Lk�����`R<M	6�<R*�z�7��x���jM�iv�my�?���,�nJ{��Mk��|��0{�����4@�@M�8�������[/��Q_�~-�c�ӄ���OeB<�Y)�O��ǉ%��q�L$�)7�)�hm`��Hz�
�Z��#�/�g�zc�{=�B5k`Pky�ѡ i\߉8�t<��0 6|�G����s�X���E:�$8n//��Z�A��;�� $��Q�؊t�� �Y.�bk71��K��s$��#�s�A������W0����by���vS���.P�ό��~ rK�$RJ����C��e��\:�d��W-�r� $7��R��,��(.���re4�:.N�g��g� ΍��{����!޾�99��($f�Xl?j�Z�LR�t�m5�2��gk�ɗ?g��DJ�1 �Km�ȅ��j=.
�C�$�Q���z��m�C��b�a���D���T��)9�ڇ���Aޢȩ���� �b��B�s�髬G#>��ֽb-��1_�)fw��"�G���K7�< 5݊�-��6K/A���.�*�kTK2t�������K��W��Q^�@D;�L744d�dך���� {�B�$RH]�5���Q�cw�k1wP/��}̦l��Y7��� �!���.wAaasd��~�܉���5���Z�p19܄�������ȟ���Q�xc�����Ea�A!����-��3��r:2�}:B�O�p�qz� `\�Gр���TTk�Q|�N���E�e��j��}�#x���� =s�q�R2���	��!��w�:����#�y���Km��	;�/�a e�l��J�-�6[w̖�#�.�H�Bb̫^��gO��Y�PX�o����<�dl�������igC��` ���6�Y���"��{�7dz�K�GtN�ⰦR �w�R.�-<68s+fC��Bv����Q(@��_�re����}�kG{-^#μ�����9�Ug��y��I����B�����6���.@}��R�J����&��L��T�$�Te3o?����H�c�7�ˎ�v��թ���ї��кHd�FM(�� N:���_T΁���l_~�(�8�\KW"��H���D����l{:&S��pǾY�8���xq�}�P ��i�E1Щw���,��
��O�H�D��k1��V�`JN[�ً?�t�9T B�.�4=̃u�e~�G��u��	��'�Q�F�4�h�$�5��H�q���	��%�Z��g���u	V$�o�i�ȶ������ɔm`�D�����)��Пѕm���H���t2 �q����r�N��K�������=�BI�E�"�Ͳ�ȨPU�yՠ�i$RN��	@���j��h�yS9��~�b-�x��}���Z�J�ċ�ۦ��K��/N�3M/_��,�,X��',�dh�͏�}���[�@m���\�a�Sah�����{q���ĜQ���]��+�	 ��H��E����H+P��L|d$`��keJ��P�F�s�`ˇ�-��gP��t����\���R�>d:�9U ���Y����ר�N*�������A3���� _Aw+��0�FE�Ww1�r-���)է��2�E�M�/Lrn/�I� D�~���d�"+�ާ_���Қ�w��
A+��i�wI4Bd*��e�?^01���!�B?���P���X�B�� \����#�&��4qh�������,Yy��/qQ����k#o���[l��=�c������zY@��W��=b��~��b�`�L���'���v*\��C,X��-$�!!�/����?��K�wp� �R�kj"l����-ҹ7�f�A�(�%�#���6	_^��5��f�k��ɴ��s]�	�%�_�;��Ҍ�� �1��:s!�Ν;άe&Y�e��L����$����������9'b|���+�}�)	��ሺ8T��rnn��d�
<��)�e�h��|�	��G�}c?����]���Z�<��ZZ����\)5;��\��K�%$�4�����\���i�(`� �ce���0\)�I� ����?�gs�Y/��T?��j�F+EQn�۵�Ҏ�E��ac�g�Y#��b���Zkw�_/]��*
h���S� l�Dأ�<v��Nv`Kd�_W%��y���f�d?c�\]YI� #�^	����-K�av��K�B��p��-�_������-X�/Tm	� �)`�|66�&^@�����,T����G��2/���{�����ۥ3��W������Ȋ��[$�w�#s:���Z٨(�7�P"��w�~�n���A]�BY��sB��F��럺%{�h�P���p!��!��v�����8EY��nd[�.�
�z�4`���HDa���fw��e�L�* :�L5�f/���"2�� M��H�o@��D�,=�Ӫ���\���*y+u�p�v�N���CM�q%*���v�E~��M:�"A�b�����@� Ѹ����N�� Ye���"���^
������VL��� ��`K؎�a�K%kNo-���/�����Rs�~�o�v�����3-R�}����0��#��r�i���e�i$��k8����=;<����خ��W+V��>Cd�O�>���\i%ӵ��h��Adk�b>zע���"(��5��T�u��d�f�)~}F4C�#��)"���FsY+$Ҽ˩Э����Ъ�����e5��A�U��'�u�VCj�8��$���[99h U�J�A�,3��0���Z�M��m9�\K�L�]e ��]M7a�?��(J�c<`w�s��T+O�s�^XMi��g��?�S���-��~du��V�$�@�[�9 B�������^��%���H΄���<o��֒,+���~���J�L�U�ݻT,��+���؞��G*����Yv�]ߡ��ɲ�~�tځ���[s��5�j�	73�{�-i�(���P>�[�KMS_K?ӴWѥ�k��矠!��I�Ǳ�7J��8me:���pv
A!��]��2�	M--��C�nB�3K�>/Sai@��=מB��J��I$I�]����9�I�6qi�a��m\�_y]X*yrxC�?�T�$0ӄ��O%m���fAC����G�@Vo�a��gO6�e�Т7�8S)j�|��0��,>�~ z�c��r��k���ɰG�@UHA�b�=���OF�2��=��H7&�Z�"2�$�q�]� �G@0MJ7���]<~�7�teF��P��d.C�Lߘd������+��L����w%X��`�tg���}����L� �n��y��
�
�5���WVn�/����tӗ0O6S�O��9r���w�O���u����A~�2X�j�Gi��Z�(o��7_���D�����w��H��(�$���`��	�6U%�lR��[��T�;�k��-P盇!S��Hm��Y�W�1k�?�M��n�
ǁ}9�6�q)���+MM��2�;õ�y:
v��7� _q�k�'}V�c��,�kV:���]�]�P�_ld��ڽ�5�*6\�d�A�ö�(�"LL��9�F���-�Λ�(�f4�F`�e��^�Q:v/��trm�Y��`�	ɓ���d?���x��S���ט874	�5�]Q�i	��N�A-�R��*����t1a�7]Ry���yo��b�V����Q�1m���i��"B��A��ݾg�u�Ud��	�����pDc���!@�Hn^��_$��<��&��p"��)��(�����5VGZ�I�����A
}gT'����F��11��ͧk�m�N�׫F��4��I`
(&�0?X�Y��`-F�7���?3��n��(���< %�X�Qp�6���mM
܎�D�c�(lCo�}&���9c�ȍĆ�0�Ȩ�='%�eO�{����wf�z��y���î�j�F��&o��x�Z�zMP�6��'��[�w�t�(�BB@2��:�A0�v>;4)�8�H�I�8K�Ȉ�Ol�Ě���:��P�+��Z;$r�K�y��{����8l�6z���cn�~�{5+��`��'`���yo�	\��;\ó�"|��M���sd\�%d�;��~=�L{6eᰋ�x�4��,�����k�DH"�<iR�!�7Nb��;�x�5�s����a��Du��Y�Y&�1d���v����1ZE^��6�;���*��7�}�)v� �?�K1�yw��8gr������n��b_�֠���V��!�{1�ʊ��X��M~0�&˞� �S�;^��t
:O�{	�c�nƍå�y��/qLm< �� D��ôgh;m���V�����g����Z�"���v�ç�eN��D�n�8/�T�/��]K�/���x*� q�C��&:")����!�M�@y}?������G�ث{]�c���H�l�����ɵ������ɈL�)�t�C�+c���.5j��|z\)`���OC������c���+��C��?J�)ʌ�@���]�3�UΓ���o/�O���%���l�E�Ѷp)�,�ɜ��|�_W���'cX�YD�;eG~��Ću�0����0YѺK�s����Ǖ��MesU�QzD\�B��o����	}��1`�;���ՀCBҬw�����U(�ΐڣ�����?��Wǩ�Wkf�[<���C""��@���VN���h�����= ID`x��W�6�8c��{��Բ�;�7�=����LV��&y9��҉
D��YUl�����h~f�jg���~�sU�n�5� "{�a$67Ț�����uU ���7�E��;o'�̹����_}x������e�D�_2G��S���y�÷�[��>����`��n����rN��
w9C�}��9(vH�t�,��V�>NPX*Y� 	��W����XZ=t8�*\=���y�4�G�fu���e� ���5*�Z�Y�tl#\��5d�+Q��/����V��l�`ĸ�{�7lt]I��RU�f~�nտ<��0!Q��<��x�NF��� �ͱW����]�=��k5-������;����'��|L�(�m��p��j�^'������/���Z5Q Y�����=��1�/ꞃ�����{/���s�Ĭ���VDs-������{OZ� �T �vV���2��o�C���6.jj����%�t������XJ)�	�q����?�4����2�$iv�x���X�FxxlN|;M����������F2f�� \E�A���j�-�DI-�^�B��A�����	h*�Y�lx��A��	]�d7����g|�8Ju��rƩ{K"f[���TF���'	�HƓ Ti"�D �,�##���,|���ԛoO����و7-D��&�U���l`�'tt�y��\��A�*�$��]{5�� ���5h��	�"u����"?[��: !D���3�����@�Y)JhU2Su��� J"YHH�g�뷙^��Ei�U\u�F��B�>��ް��F��������j�1P�ғ�ّ�@/ʾ�g�b��>���bN<-
�����e;���S��Mi�,P��8�ͧ��n��ڮ��"Z�IxC�2.;���F��s�Sp�ǹ�i�k��'���y	�3��X�C���W�
���h��3��g��B���s��'슨Eٝ��g�W�T��ˉ"��~���L�,l		���#Z��uIS�Ep�O�������WeP��֤�����F�C�ܬՙ�]*�����e;�껡|G��w�%�S�w�Ş��pǏ��*�1�S�U;���(�����*HT�W5��+h��:�/u��D �M�[���T.A������pϭ�/n��{0(i+zx�>�[�������$��u3�}�q�XT�k4��M}�(�������4{GJ�X���a~o�n�ĎE�3�-�8Ne�j�*�_mg����>p���>(��L3|x-��f`����p!p��+'���N��x�{�M�$�=�~JC��^��4x�l'�/Ϧ^�eԎ���+(1��YQsγ�9�d 9v�*Ψ�A�n�P���8!�1���H����o�P{"�3����<э����޹�7-
a�^����\�;��DJ����E�B�G����;O
��w��FJ,,�~pdR�x�=O�����[� A�T�M�NlB�4e<�S���k�y0�#��+=3F ��)}���Ϛ�a)sNm_�lڑ`�Z�x�-`�/9� �[��l"׫���d��L�Լ��L�U�#�^��5��L��J9��
h'�iij�Ĺݣ$���q��tT���hJ�͡�n�.��ەq�5�Du���Qʭ����ak)�b�
5�y������*�5ۿ�����$Q�c0�P�M���^��.9�r^�����h7DLL,�����=�U�
E)?�i(!g�+p�UF:�oZ���Zp	����7�JˍRhk,T2��D	�mkk� ��oy���������E�c}���aC�d�&���aZ�q1%Эzgؗ���.+�ܩޙ2�{|�����}+Ľ�� Ǯz��q�;`��������zRB%���R�ͯ�r�=���9R�- �^a�o~�j��)͠E&F�/�f>�%�> N܅�_c4��B�"�cajg����-��ph�FʜR�_8�֋��+�:���ޝ�+��FY���qnY|�����=�V�)���;ĳ��+�����_�H/;�,	�￧4����ؿ���D�T�+n�=�W+���F
����=?�d�S<ـ�Fuv�"������Hq@�>g&��^o�Z&�/?���f�%'�Uٱ�e7TԚx?Kb;�+,�j'
����p=��eN�d<�w �S�E���$�Tn��6���J� {R.��Cvˢ�T��=��JXJ�J)u�u*����؛7@ϔ���LKB�J4�Ji?�.'���<`��-�S:j�Q��;NL�ƹ	W��s��WM)eyEC���3��W#y�t�cz�*x��6߃=��Cc�MD���5W�?���8[J�*�@K�˾���0C��Vh�x^��[�s�����p�	"��D�I���K�Q!�s��P6o�w[����3��)./�ͩI�~��cH[ʕ+V	R�>�xjݩ͊��
���dq������;����3t����d���v���8U�ک>�/���`����,�~�?�}������P�	 e$6lo�o	��io��K��H* e&d8R��f#�l�׺d5yn֙�߿��j����U'
���DW6,����SKU�m�'�4��U�`jF{�٬�#ǮJŶZ2KT�(A���r_��KB������o<������V�y$�-�FE@�.<�-��撐���r�Ox��aWZ��&��Gt��L���!U{��t�h����P p��ȡp���_S���#�<��X��e�ƩC�Cf���N8���ܕ3�y����o����a(<<�`5�1������j��>�A��j.�[U?�Ҫ���	��[�[���
��`4
���$�Vl�[4��j�v�ߊ����7m	�D�v�(K	�̻��l�-m��y��R��4)��)�Ӫ4��]�~FW��[7�1��N�8V/�=���Fr���EwP0L�R��R���t?����?�9�Հ��xR�D9�;6"��d̼Z�O�F�&t��q�|�ʵ����Q����`�y�d�ܨ<�+�=�պ����f����.��~ԭ�(4�������z0^�>C�Y�pB��� �����!έ�H�1�{/��h�2+�WX��*
'߃��P���_��}C�Ȉe	�爝 K�ɕ��j�H��!�����/w��l=�˸��&	X��
�f�>�>��-�Ů���حP������|�G[�� ��t�D����է�aw�} E/��)o�X�н���p�9$�%|��䩃BH&�s�#��D�=\�
�5�6=o����Ha��!H{�m���'T4�6� �.�DJ�qq����(w��N��Ib!�H}���W��[��� ���e �}���[S;�b!`���?{t�PbXFa��w�2䡅~-�52�v�l���������A]�ȳ���6l���� J��yL�90��5B0G˽v��DGGFbOaOb�+d������� D��ֽwd|��n�����`2���e��8�!�����T\N<��BZRxg�q��x>K�)_�z�P��ȼ��΋Ld��S���q�w���� ��~������U7f�Ǆ��X�{��Ndz�*|0���{�S�͕�%��+�`l�_���<ȆF͝��i���?c~?�pgaz׵4�(�ek����p(�jআ�.3��X��z&��Y1�W��^�|�'G�K��u��T�#
��.��7�8�p�hY�r��Ӟ�l��kY���}�19�o��K�F���OKK9$�I�H�ir�F�Q�Bt9����B/pl3;r���P�ذ�i:�sh��,u4Km�W5�f2���	a�ك��6MF���p,�d4�D����b�N �7$��\I��AK	͡s���%�z��@�6R�Y�'\� �ۡ�� ��Nף�F�,S�ᇺ��H%�t�n&6�������� E�~U��k?���lt0Uw��O�A�b؉p��Z��`���� ���|c����H�[/4�g<%-$��Z��۽��� ��J��0q�\�}2��s&Y�J�����9;M�{.�Dw��8)��$���+�peҭx�UXFȕV3�����f���䡝zc��|���RqP0H����X�~o'F��G|��]���nn��jľ,9!A�������o�}�i1�,dc?�B�="�7��\��H�~�#��d�A	���~�J˝�͉7Y�/��98W0�����c_y����~�{�Me�s)F�Nw|�=+��u͉��>��m��(^IN�=��U��D��F07%�V&Z?{,�ަ�"�{�}¡Ё�b��Oh2��p���j�C���m��RwښIz1�D�f��P�OB����ٜ/���s8����P^����l^ZZ����E)O]#x���`%�ñU&�+�o�uL�i�/�&5�VTS�8�D3#�L,�	Y��b@f����w�]��#I���sO�d!�����C���/��ۦ�V������~�l��gŇge�cā�{��tV<Y�V�S�w��w���LsPN#Efi���TN�]ܹL��v��f�kkKU}*mF�0��U��f�7&Ai���B%���yy#�K_��t�Nu����H��KWV�M�����	�ǭ?�$�6��_�et�A(!9���-"���ʟm;�vK��<1;胵c����!_:��
3R�q\a���d\*_�y�����M��s1�p�&��)�y�@�����`��� � }�V�ʒ��+�~,�A	�����/U9?A���n�_�)�v[���#��HB�^�Ë��_`�"��/�������2�8X��)���֑H��|O�:1�qLD��=��*��L�y����#I�&���X�=0o�J��/;R1s�Nns�fݰtc>z{� g�y�ʌ�3if�ʵi����61z�.����RM�rvN�?=��v0�:�
R�򝟨��T�LJЧ�-�a7�Z���LѨ�D4;�U14�bo�r��"���J�ce4Ɉy�P(~Q�a^�5�i�Ŕ�V<�0��ڸE�� �	�j����3�'�]�_���'��ڜYbh�ᬚ�L�lÏ���"�{)===6F�S�-p+49��>Z� �c�"�\���ߐ̜ۥ^���{��H
[þ��,�}�x��Wf\�n�X1�%�jr\�^ ��G�U
�MwG�Ś�e���Zd���t���Y��G�b�*�=��YqZ5qPkOf�v֮������:z#�{�(i�9at�E7Z%������e",�P����(i����V Q=G vo�
7�+1
�~y��U�Q|M#a�=�l�H�b�ᖞb�ɵN������b�^��Z���eO�wn���T]��#�1��%�@m�C��ʄ ��Ő�U`Im�yۣ�wj���=F��`��� W���\�.��/x8��%nt&ʪ�B�}�R���<*+�o�']I�PB�$���o������lH	����%9��.td"'b���I����ӏ�1�6-�{��9�t��`���wU����@\k�����a�ߘ����}�R��j�_�n5�߻m4=����	�
�w*hg���V��+��^��{\��\�G��lI	:�ؒI w�U�@lXf�3i�[LI�����\5�������a�}���M�/�9��R7V�QV	��$s?μۈ����!��lW���G�3�{�7����×��z�����X~��;��!3V�9�e�p����xL&��ʘ��t2&��ovt���L�Oi�2�c�*� 9����D�9ʈ&F����3U����4?pyT4
`*Ԏ>���]^i��a3�躂�������$�i�eؼ��5� 0�����sS�Y��,G����%Q��mLg�����ͽZߒHQ5�`���ȕ,K�����1F�&	V4`$2��k�}b>�c�+(E?'<�w���6�H�C&u �,P.�SheFDTT����  eS���Q�ۉKk�e�-�}���H(���v�8g��s��̲Y)�L1���~�Z?sR��*�����a (��uۓ�'}R�����OV ˞�]N��;o�/�U�7�V$ �"�I	b�1r�o��1Y�A��:0c��n�5*�hy�4���X�V1�⩵��)�iHd�Q�^�I�ߓ���̦p+���#�ޗ��Gs�#i�x�q�Y�N�r��Y�JP�vCj/��S�Kѵ� �v�8��:�x��t*팊Y�NL��mtT����wT�GN����X�o�J*'��B��R�o��_@t�Z�y�Z-��ksy�6+�G�����4ۗg(=P4W �+�W��/���BG��[viX�r	b�伿h�R?�o�T�'�rB6J�-
�@�$�:}1.��;n�)�L��sC��O���c��~��2�zKׁLw���W��ݶS�<�`���6'׊I$�b���Z����	�b�~�X��)-U^��/�xh��� �۔���"Z��=+|Yȹ���-4L^��*9Mm��6��{���W�� R٦��s�1Ȕ�P���y%F���#���R_�{���Wϼ��87#���G2��S�TDl������X|��E0Mt��}j4�n�����1��6��&�ؤ�<�g���D��矷�c�$�$�Y�Ԥ�+��Bt��)����;����cG0��_�'G")�A��%��"&��_�fv�+X}���ab�:[ؠx�D�&C%/g�dmvfr#�7�i���Ubl�*�Ք��Q�63h��O@i���sr� ?`� -��<d�٪:QvI�L1i����X�]���c�;��o��d	)�i����(O$�>n��({�����ғf�@��+G,��ʧb[o^���g/VD� �W��v�=RAW*Wp�C_��I���TU9�Ҫ���۫���;�}TK�m=�,�BSl��E�"1�"�R�	�iVBƭ�-�%��\�G:@2����q�nx�^�cG�b�\�&l��	��8��r�7;(M?�b�E�v������9�07��V1�J���uoPF�bo$Rj���J�k> �O2ި��0��ĝ����S�H��Y�Lt]���z�pmX `��D���$	�O�(	� ��m~�-jέ9��½�w))��?萇���_��h�{@�j�?�wTS[�.�9�=��5
*D@�[(
"(M��H'���(��
H	(H�^Gz�R�B	=���������q��~�x�=����lϜ{g��L�n�٘�@�/��"�O`m1O�f;Ύ���r�u������b��⽨�g����sV�]tH����_��s�
�8�wY�Q3���,�� 'n�� �'�9,Z�A-��I�
¤F-DےS�����1�}u�s��~���^Ǳ�[�����e�=�F�~y4g��[��۳@ً�>2x��Ϥ��Ҋ���7oR�,��]M�	}��Φ �|�FOR� g��U�ünۣ�����qZsk��h�Ѧ�i��X��-���%��W�1g߸��-�/p�����$����}J��8�G�.������gd�(<A���Z��As�d�X*��*`�1���[�.ݞ �B��#%nv�gά�uH�A�+3��P�k�����O'��&_���A��Km��k#�,0K@wR&�[@6�T�M5�`3�UϽ��D�/���J{HB�4�����Q��n
X K�t`^�k��5�@�t��z0&WU� ��*~�z��η��-{�H��vi%�T����A� Kp�t��8`I�:�f,L��%�3��#~z����aР�����7Dɞ��1��5�>��F�L��=�
h�4~{�·�۝�\e��]^$2��\� o��4	�k�Q �""Co\�2_F3���p97�z���*����C����/��*s��6�B� 1��lړm��5�l�0��(�>�Zl�'�韼��4��L����?���7���Z�1hQ��>����V�0(>�GK0�09������XuE)s� Pf�*�]Qq��d��B3�/:b555s@��1ϳn��8�r��3kޖ�b�20;��9N;��zވ����ϓ�+,%V����Ҋz�,�>��L���B u�dd�D�b��V���`���":�\u���M�� ���|e��b�/�]��$,�6j32tӠ����w�whvM7 ��Қ��R�K�� ���~���~��F
Itն������U���X���s�8v&b���A�H�#Yz���{Z�}�Wu�ں��U�����ҧ����)T�@2(w(,=�7��������n�	�����n� ���#p����Z�L򇒌�n�����f��E��@!&y����DZ�~�/�[ �$� �#ޒ\�;��f+'�35�K�K���`�gN�^�7��n�|B�UM o�ǩ�{E֮��a�c8�����\�`���ӹ��G�֓�������Ѝ�������7�
�V�Bu��7*4���p�hOТɫ �Y6��R����
�'�����I^dg��(C��n��~; �q��H04$D����m��
�22������i����p	��nRgg�+���휢���jv�j�k���z�Y���+����v��[�|�C!�
���Pɚ&S�i���nR׎�����Vf�2���9hw�I�m�#�=���Ô3㪐h]
�4����t. ���`�Qf$���#�`��H���Q�[r�T
9��f1�����/˰�V�r5��>��F/j�6�b1��KQ��E�'��,��95yݺ
:��n�&4�E�8��)u@W^>&�V�H�8�/��K��H�O��+ܕ@���)�[ W��k0n�kǗ�Sv~SWW�i	��uie��{=H�XX���:�_�Q�4��mCG��K�3����L24PK�Ȑ��F���kY�"Bc% ?h��.?��$� !''x*�E�x�q��e!p��&X��7���(�1���R�H��h��eZb��&�u�k���������7��US�K^ML���p5�\ݒ�U�>����S9��A�����3���a�~cZR�Ǐ *w��r����[k�m7F�pC���@����^t�W�hT?{a0�Ǧ�K�KTO[u�qp��m"�: |}@R��Ww&��.&�Fy�P2�)h�͍�"\,������#���PE��
���9��[�<�[�3�x8���3�$����j�Z�-|��w�a�k&˷��jU��hU���{h�<��	-�����$E�!�E���9������n�W���cj�"���$�o���`�c���+�'�*�,q�n���ļ�b��ǧ;d��[�)�+��Y��$G��e�r�����}T� Ց�%�ٱ�.�Pӎ�ã<�f�Vn'�Ww���W�f6]��R�4G�[6~҇�s��vôS�p�
���k�O�V�*~�I�����d�����&�#�.	�6ם*�j� ����Ama�H�eR:�R׋����<��F��
�:�?O����P�AË�T���+5c���-J`��+BI�dS�����Z��<^\8Y��٣��TMM��Tm�	�	;�d��Ŝ£��f�b���@�KPQ����$#u�\mӓ�S�<5#*T�U3��S����%	~>R�)�v����"�����e�x�
i����X��H��v�:i~�@��95j���?�f'����V��S�?̩�7�U���RA��&��El��P�{Y?َ�/?��ѭ�v��j?αRe"�2Q�f?e��(��~�A�U*��l���]��Z�VX������� �����RO�z|h���l����O����Y��N�IkG}ۓ��d�t@B�4g��tm*\�u=��O=������*�����z|CP�e����A�R����T�� ����.�kƹV�hΰ�l�,oY������Й9"��W=*@�z���9X�s*���X�)�-df�����'�/8��T]T��|��|�C�!BǏ���h�����<Ԡ>��u�\l���yúQfX�T�VT�\_� �T!C�8�c�n���>":���S1ڭA��g�����h�.#�1�H�n`�1,�g}��E{��DL������9q� ��
�s0�Q�����tY�\`T�a������OoS�Z�+zJr6xxG']���t��g�l{����UH�+L�Z������I�*.�j�V~���
��R{:��~~���#~�0�,/U
�w��-1��Q����^F���⦵�c�Z��û���=�{�6�� I/&M�;r�1���
�9�FU�&a�<;rgbD�`�1
I��}	d5è���I	��$���}� �����[�f"�|���O݈�n>��DvP��((#�1)��G�����.:�'���-X��,�h�b?�$>����:B���h����8���VE�ߡ2�����Px�45�W#�<��¢�e�6�p�PO&�8� ���;�^`��l{�jFur�P+!@����c�d�=�P����Z�3,}��h�:ի�in���Ɲъ�	��?9�JL���wjO��iL1����O8?��vrN:�9T>4�A�v`�{�^�
��%G�^�ގdo}�\��~c$�]�:���k�j:��tY?��-�zδE���i���s�j��UN�$R�U�A�h�^�0��K���[yB�.K�g0R�lfZb����}�۫7Y����+������L^�d�U�)�E>�\�ں�1r�vB�*��HeJR9�
��/� ���P�.�J[�Ti��j����0	����UV>��m?P�|�����5e���������j�(	+;B��� �S�=i�::_
��H%Q�5,6a�	�Q���ѝ���%ahȥ{;ԩ��An�c�����E	����Y�s�Y�%�Ws%�yb��ˏP�㫏W�OX��/ϗZ�焮�-��.52�ϻ�i�'��w{��-���qH]=�k���Po�G�k�l��'�Sb��\����%�& I��"���,��^�nJSY���'��c��DdA�(�,"ɐ��"��^��C7h��zW45}֍9M��Л����IG���'l��d�u�����4��]C�R�Ϣ����� ���A��$���t"�-S;����,g�SJ)�::}�4���S���m�����B6W�4��K�ȷVb���]�T��9� z1!iE�Mܼ�'��1hj�3I��j��?7�.�F���U*%>�X2 |d+	�g^��]O��O��n���s�ǓHǝی��Ʈ�R�uh�g�I	��3.?I���B�V?'���'����&&s��+d;��kx�9��w����e.�='߂�hC���+����ь�M|���)d
h�2�����/u6_詹4xI-�	k�m�s�]�_���֙T��]��g;�xs ��ޣ�����)��$ �̈XC�3V���.K}Olt{'c����\Nu}�%+�n0#f�?��T϶�̮&�6�s����N�n��,c'�/?���j�D�Y�	�ʯS�����Sོ��"W;��C]a��r)���3T�v��Lk#ߓaO�.�4��tk�u5���(Kܲ]��Qû�e,��Q�q	��N���v��nn����d9�D��\X"�v��Gt�~����X+0�>��mѴ}���Qƃ�.�]��8��'����ﱖy~��.�԰m��ڇb��P��W�9Ƭw�^[5u����SexhZ���Y�Rpj���W��Y|�%�\��(���i���.�����O;�c�s4'��߭ �W3����E(k��a#A�	�D��c޻�K�|A��Z���l�U5:�м�����F���]�f��sgk]m�Cx�H�A�M�������\�b�Y7��D/��k�����~%���z�|M���&��ߩ�Pɪ�����mC49VH�2�$P�HX� ?��=cɯ�q;��koT�<�$u���*�8����J=�؍��,p����)M4�5�~��9�h��C�"9;.,�J�:�[n,	Ȫ�%F"DO�?QcrGN������n(�'�{͓h?}%⁪[F2��y�����$a��sI$~�V[�����������[I�y��E��/M& ШR @hUBB���V�U��_�,ñ��Y}[|`#u��lI!�xϤꣾD����ѵ�1N��B߁�`7�*0b�?)��Q�?���V*Ur��o;������&��6�nx�W������~%���q�r�g����}`$�L}��^|������s��E��}�T5؞��䒗��i٣1bAەx}�E�;����c�B��I!��jHMBI	�q�$�p�݉=>�.G��O
|���9�0���wB�� |��IVRn��1q��O���(��GzSS�ߑ��\Y	'��1e��G��T�Y<3�,�E±g�����S�U�.�����VQ��?�>3=����2�O�I�\��27z/�����퇰��	�I����@tl�}�f�<Y(�$��H���C}���М'bߋ�w���p�l��H|=i!��B�O��JlFT��
���!}a��w^v,�
�����adݷJa���uy��_��yw��3��H���׮�Ɨ�,tܥ���������8��ɲ?]�SD�b��O����'����_���O�	���>���K21雔��[�G L})�_�h�C�K7-#FQ�Bydl����ձI��p���X9r�^A!i�>�&l�󱦻ڇ���[�Kuaj ������\Q�Ln�˱�uhU]��RՀ~ f���c�CjK-L$�б��L������Mu����r�y��8O�� ���0���ϭEWpy�Q�V�p�bg�o��/B��,�<��U���z���L>���P%��/<�`a(���ᾅ��L�p�*Oĸ� �ơkR����O���&Y�W���䩀P��ꌹvP�q]�BR���AgJ7����#�4�'����-	;�0ə��)z��9��f���	9��Y3�k�KmZ���jRީZ��.7���gXQ�a����u1R}}b�"�KY�U)>�_�X�u�b�����KI���d��M��uRO�Їf[khXu� ����">�%6�Ay�$���p��`�t4^������+���]kd�n�x�%6���&�?�����UT R<l�jEz��^���x߷��by�j���O$��|���ގ�	���26e��9���rΑA�_RGC�4��۽/h�U�~��E4N��$�À~�/`\���� �W�ǽ��TE~yPƯ�2��]@������W���
�����(��W]���(�����rH�����ĐT��f�����R�=|.Y��e�,�4��O���8�8)t�Ƈ����+Z[4����ꨁ?>�D$>� Ѡ^��Rkvw�q�i;_
������W^��ii	g���O,V�=��R���Nrs?y355�'��א�]^���%��%4i7W��KUX�g�dgn2ִ��x93W�
K��(��LDڟ�<�V��2�Q�
�A4j�-a�����ȗ*F]�0匈�AnJ}Ή�֔h�[���b�9io rF$�U���yRO����Zݛ	����p���mHn�,�~ms_Q�?���5��ncoxwC����4�Js^�>S���E�l��#�d1L���Uk.U䬭�Ʋ�V�Q������D�����ƿ s�	Y�hzY����
�C��;�I�0Ǔ�g��
�ދ�������_lJoj����+��5{zd���}���w�P�u��/���	�X6r��2���wW&��"z��CS��matt�� _zx<%R"L۴�nҟ/��`�K����~]��y�V�H�v��䮏�q���@����=>vQ1�J�b��"$�6���#9�N�*���9)�IP�1O���	0�wrs��/k�cs��;�]��,V�;;Re�Ml| }(o�oh�2� C��k1�c�`���K��wk5�[��^�4>j�][6��8��t:G�io�f�'�C�Ѽm��t�������3�c͡�𕀋����6ѱ:��W9n`k�p��7�HA�6*ʾw���J��4^�[@re1�������)/�U�~6��s�d�^C.X?�S� 'Yu6�{��=���^ޕ ��u�Nz��b�Pᇔ����^�{��9�����Ǿ���������kJX_$�P�����0�^[�f�pQP9�3*ok���0��FZ�N[����]�C��z����9A:�*��t��>�B!ij���x����<�N��ǎ��l>o�1��\t�����6
��?�����
?Œ:�o���[W^����װ��+'��F�%N^�Zu��k���:����P�6�P��=���K9���
^gx�[V\ҟW��^x�Ԛ�%j�;'���C���q��.����1K�*��o�'8����Ú�>�5)>��$�;��ܧ;3<+����V�2�سp.6�I���w��r;*��DL�(����]��2yz�@:�7ɍ"!���u��U7'�t]fbr�=K���!r[䑳˃��w�>�fhA���j+S�Ǒ�
Φ'[����<�Q�(�<Zc/A� ��8=��Jo�y��J�od�W��%z]ɽ8��3*�w�g͝�F;�2�d����-���t̧]�	:4�QΡ���;��R�&�
e�`��4g(�W�{�&�n�(���F+$&[�m�S�|YA*M�=f���U�D{$wN�*Q��O�Jw�+��o�N��6t	��s�N*M]�o��㩶���#���q��▬z�א�ɻ���Ճɘ>Ҳju�.a�v��me,�=��CD�\���kd�8F,�"�LQ���B4}��6�$���qV.yw��p$���T*�S���䗍mA\�{�`��gP�v��P�L��*q1cl�P����yF��-ʊZ+�sn�+����(5���<Q7��_�H+��C�2*>k�R�Vn�%�r�5U�L��W��ԦV=I_��y��|B*���l���"��Ҡ�B���
��J�>狹i���O��TGcG�v�a�on%j����z1fk���@+���Ɖe�@����������>�&����D�^k��x�3�SIPH�n���NU%��BjОd�p��\`�2�`UP.�u���jP{�]S�N!ӂ�\".N!��Y n��V����=���D$Y�>B�}�>�J3��'��/T�]�KP� M�-0��J�$��<?�K����j!��E���ڞ��^ǭ޻������A�5q����i}���^ͬ�F�|c�f�ω'��Z��w"�Y���:3��h�4m�H.)�R39Y��u�T*Te��ګ�P���T5����<�X �̃Z��$JИ�E#�㳫�����	/�x��-W
�KCJ������{�e�a�����n���y�d���<p���z����f�� �:́0������ �}�D��`���F�PԮ��L>��0D8a�\�y<g��e�h�f��?��T�%|�8�2���5�y�_�VtiB�v�r?6ʀÔ�ѿ��d\��jy���ڟ���ȭ�P6�F+�١>��.�ݥ��;V��%��������
��AC[��I�@[����¶Y�ĳ���t���:�����&]��H�T$��9+(�|muD��Df]�V�]�K����P��>d��0�[֗=�|��ZXi�P:�܊0@8�CM5�=�휎<n�A�x"�:=PT����1��ܪ��	/DfI!
UY;�K��yy��5��W�m��1�3ߑ9N���?�(">��LɫUiA���Q]p*�(T׫�S+ז'������(?���w��K� U�h~�e�.N�6�C�9��K�P���T���p�V��k���vC�|�xC-���;��׳th��K���$^�y8-U�YW��L+o�l;��.�ڪ��J ���o4N%�����7@,����q��~��H��G�s���8Q{����ar��ҭ�ϓ
{Ctdܯ�D&{
���#��/k]p����	;�r�7�@' L_T�Os*#	��K����:���4���.��=�Ჲ���J��k����Wx�e3_8���W�;Aז���m7��@�/�%} ��qA
"��	d��_��d ��m�kc��/�yyｯݬ���f{�#4��´����|_��b�Ԅ���썄6q�&��O�T_*<�{:��I�]��]�yk�
o���Q��8�=t璠��S�ow��w��w�n��~\���!��O]�#*��hq-���8�D�C�G�q|�Og6����v�����@�{�;R�x�lŃ�/L�v"d��S�.<�y���g6f�^1���;�E~A�~�%�s!�#U6^��'�˲����U:)M�u��La�fY���k,vU���:n�5�U�����H!����M6�{A�.j���ƫh�g~F��&�k�	؁����)���˽/���b������o�Y�̚����˫hm��������.9دeIn.�F��oьY�r�Q���T���K�3�2�x�-�oJ�O��)�)h(#MCK�+6j�y��O��h�0�뭱T�w~�%�Ծl_�j��8���'���a��U40�!��ܢ��5�����j��EQn^m��Ŏ�bi��`K��CCǥ[��l���)9oCt��L�L�!�v�4kxa�4ܻ����X1�(�YU<����O�
�^�s�C(JkGjX8��d� �[�)�5jiU����ߓ;�_�7�۰1	��(M�76�4mё_$u\Χ�Q�#�&��"�#��_�LY�_	x�������\+�OϿ,����G=�l�բ���@{��+��c�O t�b���涮S� [��K�L�e��|f��{b�q��$�eڀ,���p��n`���`�
�]�
`t�fփfE��!ǋ���7��ц���:t$��~�;�F��-CMSծ��X������ǊuT�_�c^��I�FXu��b}!ڽI����Yk�VFUD�Fl@��Mٰ���k����)�S��6�����>��ᯜe��i�b*�CV�/]��+Jpu�%م.�ڦ��K�Ӊa�7�M1 �L��g &
0��9�-+��S+��Q�&J��㗍����ߧ%�~m��*@�/D�a�z���"�y\�X2�Ok�fQ��7�jB4�[�s�ۚ2��k�r,��t�usJ>�34b^VuLu-�*y�c��W<tyʪ0d8�`�٫��Ĝ�2�;��{z!n��P���c��Ȩ�o}�]{䊚�h $s|`M�R��i+M�����3}���o�%���=�v�M�iŕ\�SV�>?ZL�oY`D-����k9n뙈zG�k�V4���K>ܫ:`�]����5_��=hC��s�Z�Ɣ�y��ŔX�e�Fs�	pV��0�w=�ۥ�@��Y�SE��a�I�&�i!ǜ����n]KXy>\s�ch2�Ϯ�ޡk�1WL.��5�λ����<@�uE�0�Xpۉ����Fv(,P-�@��".\�����\��ܼ��%�<�X1�W*>�C���f�'�n�߽����<P�{ ��[]&
ľ4���A�[y�XP�Lz��XJ�����fu��2�M(ׅ5�A�8J=��n��{-55����[[�����z�J��Jj5�D��+���P�dQ������h�5����"�a-	6+�"�UHTm���Y�y��u�FS����v��<�b9��=v�ѡ=љv&b�q^�I&MZ�0_ւи���XT��e{��5��aA��>� )͸����V��v��go�jD,�� pH1Z�L3�Y׼l�<@Jս.��`z�*�hJ�I�������|��E�I����`�$���w��ڡ��\<��6���}�غ���sA�'$���!=���2o�|	���95��һ!ȕёb�}��Ux!�f�e#J�}`
�O��+��"�z�N���N�θ^cb�)�|�E����Um٨�[B�"���-��))_����f_�3�漄��w�n�c�,�3�vN�x�(�-Ξ�9�"0��e����F���;7��?F�L1� �6����X�YhO K�Z3!�..LK9���g��A���[Q���|��\�#��,w�H����ۿ��ލ����m�1�}y�mÛ$&��q�q�:��8	Hҹ�j���F#T��⥜r���ue_i���8v+�vt��S��8=�U}#Pu�u0^Г��_-�=��*밼�����N�f���Р].\Oy.h ��s�P�h��W�����Eg7O!�}�>
sk��pZ��#ﵬvg�o�����htg�[�G[�|M8j�9��gby��A��������Қ�Fc8t��3/��U�(��/�X�U�5+�R�ǃ6�>�����N��ɫ�斖� �&ే&��4��@�[4���X�-r��+������Bl4c����	�X(�r|kmߴ��pZ�ޣ�zg:h7��\gem���&GGϜ��v��?9HH�n1]�dV�*�o� � @@���+�Wt9�^L[U�KB3�u�Gvyh��-4Ꮚd�T������Լ;[W�fX�(�ƣ���F�k�z5B�TFUFO"j��#�e���-��`����Y�o|]ׇ@��{����ަ�Ym��
cNIM� p�q{�ln����v�85el�RP��$ �<���u�!d�$���HO��44��o���U��+^����Z֟��;;��ywi&[��m�Kx��G��8��ӗ���R�X�9Yd8�����g竑OX%�D�Fɉ�+�.�T%pY�i�;�4�CT�U4�$|������v琔���J'���ͭ�7?�fЭ#U�x/��-Z�X�Xi$�����v��֭�Ĳ�'�"2J2,Hs��hT��|҅FJNMM�:a}��Q���� �[\\�1Z^�d���ǘ`1�! �o����'���y�I�k��j�f(�Ccs����ZG�J{�YE"i�����%B�9Y��0O�]��J�>mh���y�����`O��4��Y#��xs癱���v�C���9Rr��v:s�Wʶz�z8�N�DI��y���snD��+x!kr��&�Jkh>1���tΜ��7ă��E����өa$>���m8��f!n�����t�Rn;��@���iGb�9K�ݡ�Ϳ�%��l5l�mN
�+/^�F��rZ������4�#��}E'� ��\��&S'��n�y��lN��Z=?�����cY��X��� �IAN=	EW)�G %�BkP����P0�ۤ�u������'@�+�v�lg��*c��F{h�p�{��u/_r�a<ދ)'�X@�I�����U�����]�n�2򜎔�+{W({�N,�Dj����O���B�����H�qJ�4耓�:<@S���f����/^\���Hx �e��ܱ�'-��Íh��H�M����[Z�F�2�۾`�]f.8��m&�ݭO�i�̖>���ѓ��ޝ5�͚ͅ��ꐎ�]��A�ɓ��-�8�=;;�?������*(�/9`@�<]�Y>bٻ����=Z��� 	S�TU���!�:Kĩ�����9`�ڻ���@�oO�VK��v� ٹT�r��g���0��|�j�~v� ��a;��\���.y�,���6��?�`��:__	u�5c�D�G�}���Yt��T�$VC�r�'�F�l螬�[�nS�B)� :�!#%�+��e����� 1�.~��=-�6)z�Mk� 'X�Te=;@�a����	���˫k�x􆕫�{�n�~9����G}��<�6$,�f�	WZ[%��׹��\�^c�z�|�)��S�����x�Hm�����[$]z���Bl��p�R9��x_�sV�Ӥ��i|�]�щ�OZm�[����U�Zz�Ǐ�)�������n�*j�� ����m�R�����66�ݼ���S���Y�s1׳o�QF�s݇6����y{+����)D���s�/+P� �N������K��:^O�A}P���ꀏ�ޯ����޼�]���F��etg����GG�u_u�Qd^YY�zIC���g��� g����.l]�Fo����#����hWӸ��ǝ�;�$��?�S�\O�yVn8Ja2>PefͰ�\e)9�(˸��8�D���j�azz�
�E�-4�Jtn��Q��]��G�"g��$�?�@�s̺���?����/�xu���:8��S���|(ݥ"_�m�qR���	͸���
M��:,�v��3�QA�|���P�4�\4A�h�{�w�;�;j�]�47��.��X�e5�40NْS��U*����΄꥗q//a�XB�lx�X>�O%���|g�@��Y�\��=�{"fD��G�΀bM+�%���W�dS�ʕ�8z-��9Փm
��.mkm�~<��0�1]z�Fd��_��~s�*�#���B'����~��\::���I(W�+X@R
�jWjOAA_�RE�'5�w�*q����Țz���]�%����1M����7��[��s�[>����k�{:2ǄsH;J���"JmO�(W�'O����TSR�HsDڕ6'Q�Hך�Y�5�l.j��$����<:򮾈Nm_������O��T����0�0B:�$��[�E0���r�$�mz�pIIiR&����M���iڙ�~��W?����/ƆC���S����H��%-�)%+�
��K��U�is��ϊZ�X��q۹��&ݬCCC��w��ĳ��?wa��W�{��Z'�1����y��THGW#]��vM$�����6�Ji����
e���T��a(X���E�(�n:0��{P�����+"��g�6���@W�IU8ûg�1ѷ9:e�cf΢+�K�'�6�%"]��띢Lq������Z�H�EHx�؂�u��՛$;}թ���\A�S[>Y�[X��6����' K�t����W����Pz�P�.��T@��������+�,�R����ޑ�\�=׉=3Y�M�w%V�~�gs��Sj��O�Н��W�������X
z}�DA�V��"Q��g9�� �OǦ��s�ͣ��#>�֒���í�'b����{�}/����E�`bo>:|B���ρ�/�k�կ-.oV���SQ�ÿK�K���P�n)�It�P���ĺo<}�)IW�V;$h5m�����z)3��>�۩���C��8��s+XI�5cB�W�*U��/l������ze����k[��Eih�;n�vj���ߕ;Gm�$���-���u>���������s�~��y����p����� �8T"��!���7��?[���}��/�`��g;�9��-���Ō�|��k[;}C���O6�,\��iYJc���x-��j��������龧��U���
u��z.�8���'��p����%˜��`�{��K��-Z�y��ȇ�UznMY^G�&�yl���E�R��X�4���w�·��Α�`�A��8��fjE
t�.�}n��xFz4�������L�NE+��$�W��IC������\�j4>	�e��y�ݬԽ|�`-��1�s�d<������v1A��k��~����xJc�uYɃ�Ur"���%.8��@���90�g�D6]�*"8*Qhl#�����Xln���m�Xf�֩n�k��&���{N���ͫ3+��k&f��>B�&&E+�Sʓ�$�0�$&��(���ǯ����L
SfR�*���H��ERP3+���K�0ԇ^C�� �1'��K�#�MMM�3s���D�&=�i����?�^ЗyB���	�-*2��^]u��}���_��6c)�x���
_oŊ�T����&��X�����Sv�;|�?��W?��ϙ���_���_\��W׽�	IY�MbFb�����{�hZ��Ueܶe=��:G�C�z�d	[�Vcs�,Y;��l9?$
*�?��o�ϗ�����S�[�u�`+׹�\P�ӑ�N���b6�er_a;��#�ݺ�r��5����~��G�D��UV��6�~}��b�
n^e_%멃��4�^��z����Q���E�9� ˮ׆�Q�Ha�Q�K���:g�d���du�/e�׃\�/���[�M�C�V����;����ʾ�eԚmj��%�?Q)J��h�#��O����EM/�(%�J<��[e�ᢰ�֞�׾�*Ŕ�����d��-��?�P�f�i�6j���?�L��ea�fev{}�=������n�3R���y�[���n��kf{O���}3��;3">*D=ݶha<���_��>��9�
�l+((HZ�g�Z��j��>�m�%h�p�6Q��c}y�l׺�5AF�o,�B���#_�yv~�~H���?����vw�:F}�J�@��I��9�^���〇���$����r�٥�s�Qc�%��I����!;'~W0��UDe���ͽĆ��ӓ�QV��
�d#<�'�y3MJ�^�R���t��������}9J94�~�t��#��.��C$�3������g��nf��R�R�G��u�r��9f�F(Ok~.?�!�[oůlp~�������x|C�����Y��.�����=�uO�	������P������'�&�⻬m̈�sQJ�t���ݹ�I;}v?���?��?"�#���H�)zg���ݾpH��jS�1K ��V�P��=Hw�l6�O]1J��He��Z=2���tj���{κ�ǟ��7�v+ܔ-�BW[?��+'I���X��'�׼��>��9f��:�m�Aw|�x2�d.�`V��ĥA�យ�(�@_�%���.��,"�'�o�s�I�;0�[���1�y>�6oQ�U%���.���[�C�t�C�=�[dm��E)��-��#�*{�֖|(�L救�xUS����$�_�P8���[�;���iѩ˧'�Ӷ*ػPiB���'�-�|;�C���-�2��t�`prk��1��@�I�>�C�a~����k}�)om����v����Ob�P��דs�`\MIXw9w��6���#�K����&==�[s@w�,�U�9n0$�V\Μs�ۓ�{�b@1�[��?R�c����*u�OJ꘿��6+�El��۬�=@*W���҈����O����DY��y�Ċ��ʷ�����x�Ͱ{s����F*b�n]�����PtVn�+�9�����Ğ��S��rW���}~E�_�$+Vl{X�\w㪼�����xM��0"Xtu�b'�����z�uM��z��#V�>B��&�:)���ZZ��/<����D,�Dqf�ZJƅ���)��6C*�x�gVz�����Yԛ[������}�oH���=�A�G[/��8u�/�ۓ��ƶ�+������ ��]�|g�*y/�_K'`:�WfV����׉�a��P㇎����e�o����Q�S�R��(�

{����t��-iZny<R|�����Eov&�I�������.M<��6�n"
(i��?���9�����"G�}�[=e�8�Bt1ia�ma8�ͅ��\�F�_�v�z���ˇ�_:n#�O��S��s���Bh�[R��?m��:��o�?NH9!��Meke�ez�2�+6ce&��bg�3⳽��+�Ҍ��R�k�$/���~97��J�����߸�Е�s��L�������MGRz���~���vP�v����������)2A$�ӑ�n�ª����N5����r�����o{׸2�AŻ�I���tmy�O{�<�m-nxm*�#�,%�VUs�u1�_����>��U�V,:��=��ȱ��q,���_2<�"�V��#���#m.d3�:��Y^馻,tt�S�itt��=JV)�r�u��(=5�r>���C#L-����&߭�?�m��KܹKmh'�6,�sN�H����ҝ�m����{\T�Ua���������Gz)��u�D�
�?zq��Um#���N�kV>�g�Pm{%������%ir���b���f���C�|��J���׹�+U�m�v�6�Y�K���N�n%R�+�K��JS���Q����R�Dr,8�'ń�0��e��D�bj�*+	�&��2�������&x/�jdk����ֻU1��7ݼf6�[!�m���z]����C�����_#?��F���Iz�P�ܩ�j��C8vc���-o�EX�EU2}\6cd#"�w�%|�N�ן�������w�W��bB���޽?�;� �N�h��UYZ��������EM� ���թ�����_���AOؔQ���gO�~�wArT���MV,ݫ�W���,��(����<v�O�ɑ/K�w��)����I��E�t'��d4�"u��Q�1(�[hq��/6�ƴ��|���cbC�犍��8{_M�eդnz�L�A�a��� oL�K�.���Zn!��d3�_�(�0������_p�i0��;iӚ�!R�l�6j�༉�uH����ߗ�.���e9���u�%Ň[rž|S���%��~1Օ��{s���kf��sk��P�0aD���2_���/O�}�cYW7�z���J�(���e��K�ߑW���c7>n8��>��;}�|�G�]���;��.�[��O�������?��
�E'I�$9v)G�.��f�k�<u� �[Ju���q������Ys�VT�[H�Sf�to��i�P��/�9'Y��K��Ysi2�r���ٔ�]=rcX�.�9�)�\�L3BL��?��;���}���bAQ�bDE�"$4E�w�
� %��F���HPZ��!�"EP�z�PB�3W ��;��s�8����1₵�|��>�\s��|{f1��xx�3�|��x���3|O�iG�B�8�m���r�'�H�PG�ʱ۞�.I��Q��W�?�[+�&�Rb�`��+%�rK�x��}�_��.)ﯖ�A�9tj�̂肏�F㵂��y����1�4���O�,�J/.b�H�btuS\�\r�aolұ�q�艜�������`0U�T]R����R��N`�!���	�g�	i��jfƹHV_�6:�]~��z�3�2�g��GI nqR�#�Qg�2��C�2c�b���u
�eA
'��U4���eϸ-'|����E��+������?��/�k�?�D*c��[����ѥ���c�u=�Y���R���C�t� ��4���7$Q��J]Ӏ�6��)&a?]�d��`e�%/��.g�5fae�Dc,G+��~!A�2	-I�����r��������hJCʺYp����C��o�S��U�I�A�J C�E�^��/¨p�˅�.��u`��**P ?"z�/-2s!�y_���qE���ɶ��aݜoB��:bhQO֍�ṷ�A)�S��"����,�E4��;5�;Yr{�������dN$r��<� �%���K�i���N6d��w�}��x;�޹v�J)�Oo��q���h���~e4�P3��� 1�;PhL���F�j7�$Иk�loT�h(&�Ԥ���}O�g�ꨪ+��} ؑ���I��Q&��Oe犥���bG�mV���w4R���]꩞H��p,~;���q9����O]3^����R6���i@��<r�y��,�RW�
����:������G�{�vkn@�}8���*d�G��%t�[M4���0���xO{��<�IYf���#RE��u)�O�2��Q��o4�尿�%6�#�֭���>HJ�����
I/m����s�ט�s�1ӑ�|"D�U�˺
��(n�TF�7]��`���N�z�7i(���Sq�ֵs���X��҃���׿���{�K��K//,g�:j�1y` h��/��r4K�r�PM���m4~Fc�GISQF�㸨kB:�}�;�/@)ʛ��&fd��0����e�
�**ǷL��{+���x��8�h,,sA�=Sc;i�����#�&����J�W����#��U��0���n�y��V���N��w`x��6&��p#�i��z��<����*oi�o���_�w�_4A=������>"�^{��/vG���/���b_!����M`����+a�]��_Oz_��y��"�]�Sxy��G�������'"�Ul~3:!��+0rCc��R�N�7�r�/�T�r�&���T�괛�~��0����C�J�h�oZ�l��w�,��/���2χ�p�ع]��E��^��jcS��jR[ӄ�9�lK 6��.GT�l����v�1�N���R�g��չ̸��	 �_t�U�����,�7��Td�{�zg�#y�0���S��7�_���o�8�
���� �h�W����<弴�Y�R4kP�h����@f	D��=IIzq�ɋ#�_�P����6��2��
���W]����_��7�t�C�7�u��+�h����;�N�dN��?����@���F䩈Aޱ/���������|�f�ς��l��3B��~�ȋ!(�v�<[�D�n���AvW�/{��V�W����@C�<��y:C�3Q�2
�Q�"�So���=Gt�ܗ��2B���Z.��� T}����B����&�<��V��";��?c�4� �bW�]Ruv��Ի)��������ޓZ���IR�h"��g��^��?P���Q�ʗ�O����o�� 1���"R�_d����q�S�i�uɢ�{������N~�}�"�Z�X��W��u�Cc����{��-C��9�2ۍ�OǈK�e��}��\ 
�l�'/*ۊ�ك��w���&(G��[H�u�t���Ŧy�{�L�by��,���b��x�\�jSE*u�Rn��
��xI1������}"쾖@�U"r����A�=R0D�X��M/�$R���ݳ+ٓ 8�d[��d[j�}����#��T��^`ey�1(&!����9��2�H>Ewz��X�-M�tK����Oɇ����d��LN_p�Zv���v�nn!��ñ���^	��J �@a��Δj/�Z�V��j��8�~.]?���:�V$���)�Y3�l�a@Nk��$�r�z�a |Dws��zv��r�cs�g�
��oQ��J!3���K��+g���Q�]���oZ�[{�� ����{���M�s��|��\'~�݄v��'�Jy(����Uc��e���i����_db��B!�;sW�{�v���x����5�aU��2�}�&������Pz˩��� ����۾*oh�]{p�co��z?
�;��IC=�	��	������ {����Z7
�Fr��뤘'Lh	����fC .c�DQB�Tcm�'����'N[�LD%&���
SĔo{��k��>�9=�0u��JWJ�eI��=��z}@����Hr��Ձ
5��8��c����4�c�/,J5�A	wk�����Gd��9���� 
�Ի/�%�@q����2t��=�󏦅����f�8��Hl�&��n��.OWX���s]UV��^���9�z�z��~�F%����IK�}�d��	�P	es��/��L��d�We)\5�z�v�ґ��´�c�A��� k���<���~�W�����Ꙏ�f4�9�1]�$}��c���p�ƲT��I��|B�k�YM}�༃"r��ɀҁ�a}�""wc�7H�p�KzQV���9z?��(��joi�΍�sW�f�%,�N����j��O�I��O��������)M?D'��y�c'�ͩ�s*\ Ƹ���>�'?�t���2��H�G�$c� ()p~�N��V��`nc�R'�3��D��$��k�P��^���&&�EJ%��CH5�%�V��ӡ�E��c1Ά�٠���2=���%ÅrdJ�����3���)t\��C�Q���8 ���a�,� X~��^�@v=�
�����f���I{�}��D���o�L�\��P�#f}����9-�EG�c>����� 9ʋD�E׹�nD��3�c׻�
P��j�~�X_��sP�*��!��YU&25aL��r�eD"���~�U���鹯S3�p<���P-w� ���~�������(��Oɇ�k��U��:��C�~%�L�0������2�������N]��<�i-�9��;ya��94%]�.2 ���D���P��r�Ʊ�etN�S��q�Zɮ?�Ez6�����9�
����6��b�'2�_��������+kH���|�5!k��hV�xƧ(Ue����S9��MO�Q2wUYbV�T�2�k[�[���R�90�Ѡ0��P�~-�v�&c?�ߐ:U1<�-�8��*��$W2*ZΌ��9�
��.�k�������w��Y��M& #D�¥,��q_�^e���2c�s?\��4�?`��\$x+h��Ty��/��6�I�"��Y�5w��D]�8И���}���l��Z����}+���Uf9v%�����2ФQ��̔�0��t�:TT�,���h)[������=�y��c�� v�����QM{~�h�KLKoG�P����*ui��T��lU����ʎ'z�]�0��0J��B����Ť����ZǤ(DJy���a���)��RoM�o�w��(gP�U�6W�5bC�ث�XȰY�m��</�ܷ�:�O�z�NS���ې�Y�g�B�QPR-lK�Bi��Z'��z�=�r�3V6���V]���\Ա�C�y��!�fI���kH��>j��o�u�#�4az-	���p)�\�ei����V�5��O'����eȞ�Ъ�������.��	��������d=Lο�x��2��i��/�����	*.�������IJ�\�K	�bD��N(��N_֡��U��!+%=�f�k �m炱����B�0hԠ��Y#,{�]��4�0\ )wx�������^�Ѓ�fZrHx�*S�e�kŞ䰃,�Z�P�s1!mǷ��g�Hر��1�����PL�޺LN��R+A�R�a�� ����s��`��g�����z2���"�-�afy�bh��,�o�h�YZ��b.��]��{����x�1��k��0�3;@�n��FOf到� ��v���W�86jy�I-;�3����~����g8��������8k����+��_9��_�=���Y��|�H5��=;�n�SX�����dGt����i5�@8�Ж�ިX���g}�캈��h�R|����E��J/� y=V���aĮܵ���x�=���y:4?�T��O�����kǎ�[x��Ž1���pw_:�q6	�迓���#��]��ݗf��&��IE����^���B�aMK0D�#K���2�1�k0�ٔ�A_U4sb�U��*6��M%BW����Y�4N�.�	���m�_�b+��q_Ķ\pq|�N�Ǿ菮��z�T�.�	������ݴ&�UO��k�=�_�AEu꿪x��%�P�,s���$�p�y�E��V�0�oe�b�oPm	��v��?Έ��V����^e���:�������%��5���8sC\@�L�\�t·\v�1�|j���>ij)�`>W+���`�k�D��-S\%����M��eC�)���c�x��%���Fn���R,'���a��-�`v�#�3}��3Z\�Gk�e1�a�l����gT����>���q��n�x�

	1��{�3�{�]��9{K��	�@��
���M��O�/L���M���ύl�.E�bS�� �H���9jQKDJ�ne�U_NX�}��2����cc�����r�r1b	X^^.~2��>T���=��ʵ�\����L�ݯo�-T�DˊM��ފ�^i��&���\�Da�'A�$K2u���mֶJ��-12&&��1�7���/e`��?�>�S�e�Q�Y�U�V��%8�_z�1�����U�|T���ux7,���������j�F�WB����E�����OK�������?��?��������g�حm����g2+��8���#(�+1-�H��8>B�B�UB��2�hהPB��3����19�E�;����}E�7>yO�R;w/]�'���K��h���>�\}�v����/ND���(�r�4��R��r�N$C���T �m,|��v���R4L���фM�:�>~�����7ω�4�q��n(.�֣[���պz}���Ob��w�-g٤�c�����Xf��q��J�i������=�!�����tg�;�����A��c�l��y`�]e�R/:`\k"YT�|hX�/B̈́4�����jω���Z���m���&�ض�����[Ô��ݯ���z����ve*�'�w�^,����N,�~�{���AW~���� ������OĖܓ;Q��ЉC�.3�/�+�lj��1�ؖ2<����A%�/����Z�~A|e8�D��LWqZ-�y+���Q��/�1����Au�:_9�3�!9{�b�d����婱�@�lG��n�
��7;r;���Z�IԾGl,3�H��?�!���O�C��Y��Í�oO0hL5m��~T혐�|�5�nT��q�[�����YY��l����O��}�6���t@��O�Z���P o�����g����gr��i��ӟ�n�?���D_/ ���D���zg�Z�idzD�/�u&�/�:?��Ոsē�����hr�,q���y�c���αo�ln����fb�����;�����XqJ�L��?��`4�_�@%�_��������m?�%�
*^
lGh��[�T/��}�_-t-|��x��2ڸ(��Mb���r�����OxiA��s��M�:�G	��ߓ�
:���mL�IO�{�I�?H��tR��
�6Z�G�s�	�Lm2#aY`s^��C�6�i�Gy;����U|��γ��Y$K�����6�j�=��Or~�/�����S���%s�hFOX����c���x� U�����?��g��I1�4g,;�K��#��05�՜)�To�"B{Y��Gzs3j�ú�?��[�6�u�]�Y�9����Ũ�a?���me�]]��94�9܅F-�B_��h\_����G東/_'�i�[�x�)�rn�Mͻ�r�X�2�4�q��%�/�f�y�jH�"�Mz�
J���l������lR��_�=6�茺5i&g�LB*uCg��0�&D�hY�S��l}��VA@��D����>�ͥ@���T~s�}��މ�tx���p���q�!�R�٩7Ʉ��J�7���n�Ն��S�~��8��aR������m֬�b�~&E�����rq�g�C���}u�W�j&j�O�;��D������zr��o��H�(�|������il�;�-��}��w�D�i�X��,���W��mwB�ܜ1�9e��[�^�h��蟏$�k&
g��YD��X�"��q���18�z�@,��▓4�E���܉K��uV�T���N;-f��f��oC��IO��[>�+�a�t����U��iA�D�[E[��jh��ƣ�ԋ,/w�寐BZ����GJ�5z[��>�TR�r�i�U�>6�1E��ǳ��(���כd�:�)'a�J�V��s��jN!	��:{!h`k�x�$
��"U�m�ơh.[V��X����ΚM
:f v�����rS��6���w�-ھ�/[�/jJ.1�GJw6L�R�RUWf�T���6�����X��u��<�����T�9����XB�2�Gٙ��؅Q�U��
$� ��7����@ qY�l��/o%�D�P����X~�Dw��h��w}"(�q�\ջ+n��-HǋhLfxv $?��Й���D����1��Fev���.L̀��A�,�!�����=>,b��AO�Z:c��}�M�^��1+�U�ՙ[�RE��g��ތ�~vS��[��T���7J��l��.���fqȷ�2-*�iRC�{�i�1�������8��<��Д+_�v�E'!�A,���e���ȎL`�J�\���5f�¯����/t1�?�R_+��+"�2�7�s`�ki��}u�.��.��K�b>+e|���&}[�h����V@�א�p՜�	����.x��z����i��&_��\�n =��.Q¯�1�OCe6�}6]l�A����ͨ<�d��1�p���bS��u��	;�kS����������������W�1���mX#'�`�r,����Q!Ĉ	{�W��Ȱ��.�)�$ljz�˗��y��S��l���1{(a|╰f��w����ܛ�3�p���~l(�rK��)��N�l�mձ�K������R�h�3�`��a�����U�rub��0�!�O�+%��}�̊.ݠ��B��[�(�F��(Lz/�n��T��2'���Phk��$ ˽����!�n�ܯ5"Ν�fLpXq$º͙�ax��v��ծ�~�|�V�9òc��'?(��
ԭ̱�*�8N���6l)�=9�B�0>=9�3H�V�R?�z�%�K5s$7΃�I�B�fj���V�N=���L,raAӼ�
�x�a#S��
����q�Hi��Չ���߀p�Kq��#?��vm��LX]���=ej��bi�l�N8l�ϕ}�q|8&|[�?H�Ŧ�G�N=#�A�Y,�OK�u�x��ᤸa*���?�"�mH<�m�s$�)��9�ߑE7�����B�Y��S>��?ĝn�-��A|�O��r�>!�dN�L��?�^�<�t�#m�G~(\�+�E�x<�~.�<{Ǳ)��K��O :?T"}D���p�\��y�q�T�o���ʛ�ג����shu�W�'U�s������5K��<h�}[sL¸T���hB�Z(���N�D��Q���T�N
hξs��s���/��;�&��^�}�Z�a���3̨�o��=�L�
�{ç�*���۱Ŗ<�u�����%�MTM�Z=�g�4�!W�P�)S"z��H�{^ϓg���1,ŚI��'ɩeia���nB�v�-_�<��T;* �}�#�M���͒ח�}�?�Iռn& ��>����4P.4��h��@I�![w��9���^�`��_CD�uޖ�~��70� ��!&�2���k��}!�~�I>C��᛫��gyv�D��I�q����m���[y�ՒϮ.f��5ka9�,%��t���x��(0��C�*+",��=����0CW� "Ӫ��ݮ�����Ge�Y���q|��g�A=\v6݋���N��<cm�RۺN�ٳ��)C�pͺAݞ ���[�V���S��N�!�~����e��_�a����>���z`�WW�+
d�C��!���~����%��� f�VG�(�Wˤ$�/
O�2.f���V��W��}�k�Eԏ���UgD:n@��a��~:���6h�ϯk�GuZ╎��t5�T,Tcy��������Q���m����=k��4��9q�*3�_H��q��c;��٦��,m����(�
�|,s���e�
����2��X8�0H��Ɉ�KHƦd ��jvSVU�G~���CZ��eXE���@U�{ٔԫdP��<��~}
��k�V�釟����d�3�|{��{
��?��x��ti�o�l9��3{����̏���R��vp�,�Cy��#�\��{���6�e&ˇN}�ed�춭t��.��u�6�K�N�4 ^�*fTw���U��u�詚��)�*���<�s�����F5Mҵ�܈ j�-;�h��~	�OR۔T�)'������Q�khL����"#7M�u���Hi�ڹ'c��=+:?��z����U��Po����.)��ʵ3�<�<j;=%�Z���+�P8hFup˼<o*1��$�q�*plUPFZf4M���j�,q ��26�b�+�@�a��[~ئ�c�m�U�R_?tt������c��!LB��9h�D��je.�!����%���-����M�����{��t\��V3�j�S#{�'�v�5G�<�> ��u�%=K'N@�o��^�_��&�9�>҅R���x���B�js�04���O��@qҫ��Ɠ���J����7��Ep����	��HY�\�j��Wq�^��_�����|�ٜEZGvu�^�yڻ=���4���Z��[Ъ�w������D�� e᱊�=%N~)���zji,(�~�N�t.4�G��M4����|�\8�$�VR*�f$9LX���:�4�0���Dn���R~���B{_��̰�� 8Pc������:fͣtU��NUULps��(�|��w�`��[|�!%���~��aA�p
���΋nE��[l t�cU��׹�;��ih+�y�@�����N��[~qPϥeY≰��
�8�Yc�$&�؜�9�kj�2�K�O�SP?���T��C��'P;�sD�1G�n�QiIr+�cU.�B.,'���uU����nb�\\Z*r�� �Oi���
h��0[���Pă���WI)����F�4`�n���L��Oƿ}�t#!ͧц��}l!����Ufc����^m_��Q�����@���� D[�N����#A4M�-RO�Y��7`yO��D��(���6�-�F���HbR��|b����
��+��g �,K��:8p}����7?��0��]˩MGa&cu��Ft(�j�䇞������qL�ӝ�t�ya���d��V�`lh����Vg/=�́��$(���= ���2X�k�o�)P6��ޠ�7i�-�+>�ϧ��a��o�.�����Y�i�����R�U�Olŵ�N@�kG���0Az�^(����XE���?��zS~+v*�j()&e�(�A�����nn!�>��j*)0#�s������a7�x� ������̉����[��eC�I�xq�T-SIY�崩c������;fR����sm>۔H_zo��_`u@_D������Ƣyކ6�QfH��޸��TS��|#띺ܹjt[~�o�Y�R
�Nu
a�Tj�� ����K.q�w�&��粼(��p�N��O'� ��Le�'˾ڔ���eϦe[��������#ݓ��Y�t�UieP�t~�'_�B�B�S������	x}z��)�U�8i�Nd(h΀
1������sQ3U/��"ʽ�L^�d�7�K��(����˄���&#�� 7��m�g=ס6��^*����`>��
��V�9�̷���&/ٿ�![��[��w�!:	���t��ƚi5I\4�E�9����d�n���$�'�ʗ:Y�bퟺ1�l��5�y��ħl���˻4�JW!UNZm�mu�?�� �(�JV�Rp8�#'\
��,�6��Hf�SF���x��]Cg�����R��*hIjK�Z�̰N�W�@�I�z̷�H�b�⍟�V	+Q�-�e/��U��g�������;�H'��e^ӱa� �i uK�_�~�B�H�y4��{�y��� ?�q./�u�_[e#�R�#`:�E�|�a+�~^�R�@4���� �D�=:�WPc�Ҕ���ضP�y�TA��n�h�S���a�qu�t˝�*m7��N�\:䷥d���+J�C�Pa�*\I:tM��.9�y��r��ko��	iG�^�7�w�N"�ԏ����}f��j�Y,4Pz�3`��A/��m�
����ގ�� ubL摫OK�q�dq�J�CT�/$玲����Mb�g���
͡�YR��/���/mTd`7�n��d��xP�)Q�W���ؐ�wo�����9ض�\ ���wS�:Xji%ᤲ�X��-C��wÌ�:�e��U(߁����%�?��#�y�iׅB�� G�Β��|�`��T�TGR2�{��j�-���`�h����:��ȧ�.���C������P�˗�׍���}�~��xt|l�Y�9���c�!L�cIs�Ҳ0�;�[��2���4��������gQ�����s��1G���D��>MR��۱9LS��`����f�|���	�Lʓ�UG;��;@�q^�4����w�|��+I�.�Ѧ`'�ZͰ�g���$@,PXn#�-��蠖H��	b�:�[H�}��^���pQ6��������G9�w�*�`{3yh��^+�8)����l�.����/�a)\�]�*�1���'��h�i�A�SM�X� �vt�@�%�k)fa�Fux�kt"1?1�u��pV��Η'���Ql{�Vڷ6^�&�B�[����g����+�F��}w'���	e��*�~ЌY�5������z�Wf1�uy�E��s���?��6���XB:���  �uA+���7�����+G�T��a�J�+69��y���!*�ѽ���I�J�Of�a(�\"�͡�&q��F�p��>}�jf�H���|�18U��DfbOl���1�(A�H�����V69�G�����k9���?�mh3����~�� �R�zM��	� x�k ����@����GuѺO�D2t��m�8k�t��mщT�Ԏ,�p����5ӎ�<�mX�ba��6tT`��J$r�v7M�(��m����"�:�����u�a�2��{�tSt�|"6����EM���9�-s�3��lE�+����P�],��=��@�%��e0Q:�~gށVtr�i_�IKmQ�̪�C���OȌ6"o������X�uF�zeB\N��G�D#�c�V�|�S�C��m�'��P�'���7��u�C�2T]�)�~yX�R��ab�x#A�Y�؄�����Ne���Z�.����8��?М~�m�8�?���:�їc\�r���\V
�إ��	�5�^���m\v÷#4�_	�Eԍ5	�Z`i9�G�Q�I����t�o��d\�i�
k�C�����b��M�iuI7@���8?�*g)�<u�����6�p��G���<=�� 4xg�ywM5��%7��4ԋ�1�(���)tnO%8�d���d�l`<�d�4��!�;"-e^bh�:W�s��۔3�h�e.�L���������!��LN�*u_r�oR#����z�9  �(��r����<���Dv"��)k���~ꑺ6����PE;�Qr����q��L!�ۏ���Ay���H��A_�)��&�l��w����I�M'���PQ��f��\�XN@o[��<�
��.����"JіD����bX��:�`}�n�+����.wծ����"I��m�0��®pZ`�u'�8ծ�i%1�+�[�'�@-C�Z�����e<�T8�1E����X�����]��u�4�P"�!M��k�����{�n�]f�	��ֱn��ׯ�Y��"�*�>���6Ƈ��D >x:�tbLї&����A�8>���gh��vf$�j�����itYQ�ϙC꼶�F?�zkZu�r��Nӳak��k��,����d����v�h�"���{u��bϽ��������Q���!�����Yi�)����~�l(�ӛP�[�"��[lr�Cy/�F�+ؤ��6�sJ���;vN�Ilz�ne����U����[�	�[V��)��#�ޛ�ei}NQ���B���\"m}zNw���`�Ƥˢ��ո����>{w�/�� �,�J��]����C6vLUp�p��A�z��ą����^[T]F���ͣ�S�M7J+��T
+3������p���u�t[	���|agjG�|Lh��{С��xoa]��"�J�Do������;9�<۽]󳶞�Kȡ;;���.��z�ۄm������UO�DR���[_p��\��Z��љ�3c�*S>�XyjtU�É�Z!��|sɃЯ��<�1#����L%�Q���Ȧ�iR<�@n��uwJ���V��t7�dt}�v'�(u���3���;ەߘ���LUn1宧�����26����W��Q��"�s2���x�׈�	qƽ���e\������7������l���;}T���,L�_���ᰲՊv�<���u��u���JHZ���S�Q������."�]�FK}Ɯ���P�C�%��35�V��#�(Ƕ�ve��ں����%j�T��o�������\�C���$Of���=�2Bݠ���PO#)�z8i���D������X��Z�&$c�������V�����6�,옍�0��U
8�57ֳ��?��N�� +�-��	��4��R��l����`�/(�mU��6/"	d~�ݾ%��rw�왱6@ҫ���L-���B�͔�jM�F��ׄ�˼�ݎ�'��]{IR�5�xam�Ys�4���͢j���3H2� S�6���p��[n�J�B���sl{`�6�9r�J�-11��EҚ/\\q�1�u���C?{��pS
�xr��7_-����dn.	Ҙ���U�8/�:�l'��d��U�Fw�er��J���?��يl��P&}b	��YX%i���fz�,�������.������Y3�sU�%�>�j7��Hh5W~'6�)��Kuh
�N&�����{/M������C�2�"����PE#��=i(����b�d��W�Z��/kG���
�9+9�a���H/�����*Z@d�즐�v╽�PDy��/�a��5s���m7(&)�!SAz��wy/_����{g�=�	\X��e5�xA~�Qw�S�����O��p��`�����B#oV�V��R-����(3�읜��EE�{+�z��Ā|��k]WT.��ӧ��k,ct@b~���g�WPA���m��/ވ�����Z�T����mb�h�lx��3�:��*v���6"�s&
�bǆ�C��Y����f��}��F(�v��v���{����,�������|�SKcoίz_o"G>I���5��хNc�Cw��0	�bAm՟_�����$h�[Fr��{�MB�i�oVlͷ#,p��w#�h,���<c���H���x��M�}���]~�z~�e��>�@��;�>&3�k�u��T*f�bt�^�#�xv��b����bE~z<�O�©e��"���Y[oM�F~��˸�j2VY��N�bMx��l�Wmkh�Dm���p���� ��!��{a4僥}� g��Pg��j��)^�b32�a��w�t��M�03q',HLL	H�\[b:�h(��zR\���;}LS1�b�Cp�U��\Ut�bݤ�B��EU��:͖�kQ������5�e
����?`���S����8(�<BV����C���ǝ�z�d�5���&_��	�t|4�łH���f�Ά&^��k���U"~� Շ���X�ʅc��i���Z���i��Z�R�\�f�g�]�>��O�~0hEsg�ě\ߦ��S��Z����A�]fD��h��������o�����d|ǔT1���H�7p���b^����_���$��SS�$;��,���v��ɤ��G/s�=;��t���,�<zVP>=�J��Z~������1{�yܻ�4�VyGւ�|"�J��lqo�� ���.��Ü'�Տ�ֹ����]�h�i�������4{�Dp8�Z�<]b���.{y��1j�����F(��T4O�d�3u���s���%w/��L��ֳ����[u�\x�����m��*���C�pYp4��gB��](�B�?�t��C�y5%6���0��чt���a����db�QgT<F-�쮍58ii[�&����o��H?;ĪE$����TX�73����l��ɴ�W�V쁪�����O�|����:�6j#�V����4�Q��9�{�j%S��Vl܉=�(��j_|�x�VO�P�G�feK�_MGy�q\��3o�.���"����Q[��j+q�W���ZU�S�	�^��M�"ի��{�T�c�3��������	sKn��%�BP����+{.�	��4�ύD�L�<���CΕ`x��^����Jr�};��reIƄwO@��{6�v�R�G���-��>���*6#��u�c�=��c {�̈Ǎ=���}u��Խ�z�����tͭy���t�׌�ߒ{�T����,��kW�����T���C�aIIg�Z��s�$[X�b��tv*+�qB"M<ͯ����V,�OTfK~ݻޟ��z��N�ŊE�CJpe��(�̱�/HL�O������O'�[/.��҆���+h���nqOav�#a��rۍo�zgg�MMz<Ή������e�(w���4���UT$�Z9�nʾ�C�Gk��:*vRC�/��n�?aR=���>s�����1pS������ݕ��<�g������;	�rm��%,���K*	���J��mX*�w�Rǂ^�q�����R޸�{�<EH�H�����7�[s;Kh�tW�?q�O��C��'G�W���Sy�t�k�z>lq�A����Yk����,�]�)�\�1��D���z4�%N�$���m�m�$�A���x<8��m�Ɍ�ʔ	14�i�3���?��pp+w��碌@��X��t��\�{$��Q���wf���obΥJ�=Z�z�)�!�d���ѶB3C9��g�#ḡog��cd_S>��'��w���n��dvv� C�m��%=@���R5X%�ٕ����=9�E�ШV(��=�� ����+g�Sc�b��+��.���-a�x{y��.��ɟ�:��Qm�'r�#5=+�V��l�H�(���@�ѮԨ%��m�b���ߥf��W	䳦W64
eu,��Us�7/rsSc�WGƍ�����,8_4.�p��G�%҆��~��9��6>��,R %`���]N�V�F��HA`��Q�8��~s���ߝk۵�Ru��A��k���q1N����5ImX$hv\��uD��ԑV�_�2a�ۺ�I�Iw�32���L���x3��H6��������2ȣ[c���~ye���`Hp7󺣜q- =Ȓ9>s�zH�t6~&E˹.�%��Ҩ/c�U�E5V^D�a��u���N�K�7�Y������3�w9þ��ߔ�u���C���2w�c���]�fK�J��Dk�oV���n�i��v����g�I�춳��H[����<����2h��>����*_��r!��˜=�}��k���?�Lx>?r1w�A=�*f�]�i��+���?��Z�j-=�[��6[K�s�ۿ�'*$�{��J4���T�Hx�i��写��v;xs�G��3P�9l����+��C!���^G+�y��Q��!�2yZj0�M{��$�==Á� ��߁�T�&���|��kC����'��S����Tڸ��"^zjB��@��i�u u�$En5U���� "Pu2-o=��������g�j��M��*[�6���l`�Qj� �Cc��^��/�昑(�v��S�d2Q�U�wa���ϿjP�i�`��HÇ֍j��Q�G��fY�zZ�R�(-3��8�xX���tQ��B��k�{�U%�iq�7z��Bh��g
���o������k= �u�Qc��S��4�� �c�0AN�5W�� Yz5�g�T5h$���h4bq�d���1Z��%z��i.c�:�uC&���Dzz$�E�`�߾g���4�?�l��w�]�o�@���/fkeU�{�yL��['G�5`ԅBCӞ3�8a��,W��9�$0�W^	|3���E�7���8ػmX�����[��ڰ��'��e@@ ������3�,gf�dV[k�HQq���y��� �[g�A�l�XU����6�:��_�Pb�3��k�g��[���D��p��o�NlPU<ن��](;g̾a�g`<Ei,q��?c�� Y�م�V�@^e
Xy��Z* WZT�4�[�!~����O S({�po2�}��bD0��J��CO��Ae�laV�"�so�JBl��U"�%��b�-+�6%�/��j�\d�ӳ���t��3�����_����D��� �Yx�0˝��]	�R���m��R���᠒-��������w���V��yk��-o���Ox���ڊ��a��QU�E�'��oC(��v����RjB�v�?���#��x'�Wa�\mљ���e ,W1X�Y.彏�Y��I�f��XE��͞�tW��RgU]
*���|o����w��N��j�g�-�H�:���'���=�_W�MX�i��sת�ً1VQ\c).��K���[��rwm��_\�k�[D����$~}�������H}�3+�K't>�O��a=l������.=UyA�	Ya��tSt�R��Y�;W���[4�&ZՠǛ��)�	���cr�@ݻ?ݑ���ͯiX����$���=Y
���^�q�]c�����>7v�����y�Q�J7�E������?S�-�^���B���]�M,m+��F�+A��[�].N����ȯwIow|(�Di��@Ttt��ґ����:�+��=P�L$�H'�!����莧h��A^�۩�yս���/횑S�w�Q�R��bc Nʘ�3���P�j�rϒ"��X��R���?�s�h
Ι�Ӯ���[}�;)����5@���6�m��2�$����r�������z��Ǳ@���.E�Ai�IEB	)I�R�F:d��iF:��r�{�{��������7�f-����>{��y�9 �-�Ij�_����a� Z�f�4͉����[#�7��P;���;��:s,R���X���l V������~O��߷�����x.�l�&��9�����=;���JBݟ�7�V]�MD�Ql�ت�Ab`�̭-�7M�R��E�e�?.��v������`��\%��$iq�&h�|0��a��u�g�ڨ��9��T4���aK��`�����cqNx{U��[�ۚ>����?���&[1zQ�����h��A��I�V����D<b��_ ���e�� �1:�_���Z/&�)�u��2�!��������{��b���,&99��'��쭿{V:Ŭd���G��z�g�P�8������b��	�8Ku����q�Q�fc�ȉVq`�7�Ȫ^�>�4a�IV��l9��ut�B��Q��v(_��q���ܼAn^`'N�S��4��4��-����ku9�Ȳ�����S�p&1��*V�����J�V�Pkh�㟡��n��hۼ*e
��#_��UW��a*����3�0�еd��"�c�q�?"��Ā�6��x�:�3���'�q��A����X�ٕ��y�Zt[�hQX`7�[��nC\S�2��ە���N?��+Z!ۊ;$$@(�w�}�`R�X�Qj�;��=(�=:v��(�Q#FGk�a(�sjx��֢������HL65�I�-j5��N���̠�%J,����ϛ6r���ѡ�%^H�6�Mq�޼���1��6���H{Nɖ@U`��"���NL&|��2{�Y����G=�c�!^�S�F�<��(*�[re🡶���,��Q�����p}u�ͳ��N
�w�~|�ڋn�j���,�j�Np�*�S��o�KY��fS���u�T6�#w��wvܷ�I��ȑ�i(��Z�<�0�'��7l^M����]]�'�z2�O9h���\��0�k#d�R������fqUR�,j����ΆoT>���I�D�ƒAm4f��$�V9)��f�j�=��A�vo�Ǘ���O���5�Z��<�\¤�&z���/F��V��h��9��	�Ye��Q7,h�VreG��  2Z⇇�
q�_�
n����#��gf���'�P���hB@㝂�Ҟ��ő�X��Mݡ*�7v{�l����dY����WQ/����ɓ	V�����"�r����w]�O���;�J���v�L].������կ�2c���X
L�ťƄ���5���u謪��@��|0��B����?�T���7��
8��#����^`}�شN�8�a��'�����B���'#E�/vuJ~���+޼���hމ�IIv������e	U๕����a�ǍU�A�#L�&j���,:�<]#Z�HB��>_���y"/����m?M�I݉s�W�d�&Z�	EA�1��^�w�[d�w/m:�o'��Jl�G��o ��T�0ub2U�ٌ�6���B�P���Pm��T��H>�����i�`�SB7�"f1��M��,b�U�+�_�\G*Z'K:Sse=�0�S��l��˸V��5:���r���C%�+������hV�iND݆Dw�K��t�C=TU�E�(�!}�8�k��@[M�=��"��"���Z��T�dr���_9̿�C)ƫ	�5�9�����x�����ɻ�gs�%��!`�IN��9 <0x�~����s�oŏuD�Bύ��:����������.%��G��K���E���=]�0�b��FU\M����dj�7�qo�I�46l��z{vVr�m�jBC��؞Í�;��h�y��̔Dv�4��L��x�wc�V����d�0dX��z� �&��s	0��{~w� +]���Ҷ��������Sd���Yԯ�����E�>o­	-���K c�}� xd �V��'L������ŷj5X�������q�yk�TV���7����=K��X�L����p�U�D��P��g�~>��8��M�q���q��?GM�$5'�?��7�?'Qd�s���Γ<!��9����9��q�������~��E�9*"�y4��y^�9��X�o�>F.֭�nӛW�p#~m=�Ճ�5ޭ�m$��ͦ|�fX*�����P
b���Q�E>��)׈7VJ|�O֟5r �R�DY-���ah�6$�V��\�9�^��0X��,!/�� [� �I�nl�t���b	@f�����*m�s
JPP�xOO�xl��@fQ�G �̻Uo9�GrN5"_��P]!�G�,�;xhKU�z0kE���*/�-��]� �Sw�^��������q�����S?���+:	�[Q[���%mL����'ۛ��W7���lp����b�_!��i��H�U_�/�1\pX91�� ��̻�����o�'�ȴ�%[Ͳ�jy\<w*9��i��릦��P��?x����()�����A�A8[��}ۨ�P�=���xf'����.���>f� �0�,�Q&�����3��`�'02z.'�b["	�q7g��&o}�sV�Z�J�JW�Qb�*:��A/�����[K���:��n���vf�sദ��q���m�&yfQ�'��/{"��_ϻQ��#�d�'�.�ʘ;��)I�|�q�8���jG��A�2C�6�xz�Ǭn�/6���Tq��l��~Y,
���`p���s<|Y��4��/��p��Q\_�9�ԠJ��~�:Ҙ"�ԗZW�����\��Rn�M?�j\f�N��@��5�i�w���hw�C\���!���rM����,9��b�>c�S���O	h���m�7tWY�΅��T���0pH��	��b�s�mA���շ�|$K���A}����R.��uK�ʀc0�J����*��
i��t4Eq�� `�4�*����kc�X��T9MM���2��w|�����6���ۨ�4��l�(E|��|�Q�p��w��ab��ˆ[o��*9iͶEg�[u��>3!�'a���T���D}� �����āo�5ޫe��:f3�\H	��?QD�ɸ���Ccկ{��<M������� ��T�n0nBh�"��~	�~gc��Т����}]��NS�C9q�����[����Bڂ�������ӛ����	dS�Nv�c�ĉ�3ZƑ����<�tt�B���f�X��=������������Nb�Y�Flt�J=0�+w��#@�h}ON���I��i�A�.N����x�|�*sT�`�i]M]*�@ᚻaú:�Ƌ赡���ޢ��b���e`��> U1yN1�	QL��}��?���<8@��J.7 ُ�r�hH�P�����H�\�͈́Q��o�xbF/ب�����>��g�=��o�mfM#Y\�n��>� �!�ie��K7�5F�߄�cJ1�K1+����9����xZ���.I$uJO-]�b�ȮȠ��ǘc�!v�3uV��4nJ������'�[Op=Z�Ԋ���(��waD��{����/�W��MN^��jQ]����}5_`���Qf��\�1�}�̼Zc�ևM��s�M5��|��ߢ�B��4�1�{L�4eE:�TT�(r�h^�KQ�0���0���F�m����l�����|z.�m�Kʞl�_��]�_��r�T�.{��H�kq��u���07�b6%�(@(��C��%��kO�R#J�}�;�67��a|���1;���)�#��&�l��6�߽�\1+�$&'{�Q�T?/c��`.�� ��"aM�2�,E��ĸ@4/��(���0��UYcn)/�f�������,�'�&��~~�{ɫ�ǹ����Z���FO�*�����􌾭��[�zs�N[�4u/<��wG$�ߗ81�9`���gh�j�Z"��i*��� �M�ʁg"��\MF�9!�N�HG	 �d�m����Q穡�'�]b������4� ��|����髟���Ft��$��
>��S'��[+�JI$�a�v�����U2���k�����nn~�KU+���I� H���h(y_`vO�� P�ؕ��V�.؄R�5<(1B��@������0��t� f�?�?�݊�r��@?����ZIh\
�$T�h�ߛ��)Q UX���)�E������T�1(���͍#U]�)t������`@$�z32��1k8�c��Gzq�Kߣ�0��b��#���ƹZ�>o9w]ii�F��8$ܞ���<�)q����5)']�y�u=A\7~�t�6[#�,�Q��v���u('A�s+)~�&j�Z@����=̇ޅ�'vtts6�шNC��Z�b�9��zu�G6��|W�f�z�hN��^ڐ�O��e�F�s97�gH%��:�?���Ǌ�i�V�TW�`��"Z�:��c�r�A�v4��,߁~�i�<�-g����lo�x���0��-:ij,��3n���#�/�G1���DPK�� K+������p0���>��a���f���^���/K��yR�
�z�2PLJ7k���2�\�MY�ԧ�1�G50��U�{����4Z���V�M/�;��&V��J��M��gݤ�S�l�t�s�xeL�C�Y>m礴;:�����fͥ3����� d��9}��w�7��坼�b]ыm����y����.V��V�&oϗru&���]��"r�w��=�gR������;���}ȃϬ�~w}��7 [$niOK-�Sբ��4ɻ1zG��]�b��7x�Ž�y��L�����G�����01S4kg���Y��/��q�N���?� 8dx+��^��-�{<���n�����oeaF�6��ۍ�7�����-Ƈ��}|?��\����n�ږ�h�YJ��x��B|$�~�ҵ�uMT��8Bީ�<���57�^yQX!jI5��pIx�j77����_�0�&��FM�XS팧,uC�:;��Lm#=��ބ"fS����s *�@aˠ���w����u_'h1�=q	sDA���� m�k}�_�pÝE�t�#��j601�F&�(I�~. ��g�9���e���z9�8�ٷ@�h'��S�	W�2�ă/e���D�%i^�����o��%K1�����?�b�� ���� Zuy�~�Ƽ>zv�=�'؎��;O������K�u�������]�p̐��z,�ѓ>�	7`Wn��b�ЧML��*���\��'���A/-N��}�	mx��V�6�)�K��ŃEr�&��l&�K���J������~��3fE󘕔x�^zT�E�-�AO�ߓ~FC?^�\R�H�����|UOr���~T�3�h��6�+�jxѽ�U�����@��8�B��6�,��3�Ɵ��v��H��xn'�JB�O�'�Ę��9%�p�����m�����#j����a��I��Q�@�
�t�[�Q��J�B�V`�Tc:i�H�k����Ȋ�Ut�]�6w��fP�6(L%x��"[��.�nxOꙡ��x�L)#z_��J@z�"��o3����y�N|=4����6#�-Y1h���-Ɖ�����S����y�$U��N8Յwd�w�����Wt!��d��7X������85���TrȦ�SC�OFurw�\/���º��j��䐊e@I]w^b�L`�J5:,b{KE�w�5��Ou���=�Ŀ�hױ[��q~)N[H���$��&mD{����'L�ml��>#�-ٝ��T�-s��&�imhV��/q���y6U���P&If�-W��y����1+�c�"��v��͇'o[<�Q�D��j X�n.�ޫ���;j���R�y\�������bo͡i<�㙙�5D�IfUý������_{��g&�8�OܺǱ����8�֣0*�m�1 �<��M6Hn{��mm�h�S�ng���3�M�臚%�MSP�y,��JV���a�kEl�E��R�s�NZ�	,��U�Tr���:e'lЉ��9Q��%
6�r����AuT_>Z��y�SmX+�k�H�#�ٗ'�t�PB��kr���9����MGG����w�f�~�����������g�'��8��x؍'l2�S�ѭ�1N�9q��輮��6���<����N��R�鈴�貨�[$��1<q���If_2�d ��z��l�I_���r�
bw��;|8�^�����m^{�
�MI|譮���tmM==+��� ���J�n]��F�Zy�ƥy@:1Mr����v)���<�ml�D��љM��^��5����B�[}�\#��,��������S�^5L6=�)�
'�ɜ'm*&\1|��ik4&�ְ;s
Us�{�������sM.TN4�?p3���>ps��vm�F�����ܓ���ֻ�X����h�(z���r�q��r?�-h:���u����e�r�h�'{�x��W�b�5bD?x�yvݕ���7����6���r��r�C�w�
} �<
�}��M�3���r{�����~�i���T��D��5�5Y��(�·ר���Ȉ���H��8�V��Ό����"T��Dc�1���2�M\B~�:��Wkir2@���zz� �^Ao���m��D�;�qX2�� ���1U[cw#��;χ��:8C�9Fl[�7t��	�N@��Z� �ߒ��y<c-�l��%��5cR�#�L���'�`��9-���8�	��

A�D�X?�9���o��z"�H��v�Y��;�r1T)����x�s������ϻ¯�c�����3�qF'����֦ㄪ	x����Hp����n�]KTo{�`��h�|Tdj�}"��|6@9;H|����r2���9�F�����5������w�����1�~� 8���~�!�Δ��h��9۽�+rz�������~���Kѽ�G���s,�e�Q@,gݝc˵̯�u0yQ �j)ʺ�mZ��3����Mg�o9����+1����O��C�����H��i쬌�,����Ha�.6i���M����W���Q
��) /']1uC�^�v:�狜����R�6L�/}5��V�걠K̩�`Ô�	�C�|�����fy�6!?��zjV���oe&���އQߋ�G�g�1�@Ϩ��[S�Lʡ�ۑf��p��V��@�b�)�RQ�fY/gn�I�[�^�c]�o��Ɉ@9�"߳^���SQT`�@��͏'-Z\�����Na�&�iV�d�t:�<�X�O���:����z�܎�c�7#e��(��D�Z�7]�^E!�(U%�k�]�����^�2k���L��݂J�~���d�N�&e4߼��e���	d��&z*�,�.;��;���K	�v��T��H� A�_���Y��m~�S����%ߢ\�w1=׫���9[P�0����_F�;�;�¯���V�fsY8hޕK_W�N��iy8����iEl���m#�	cgg`A����"���(߲��[>��~P���$����5Z��x�rDn�:�$�O#pz\�͞�=^�'v"P �,��W�?��Ǵ�o����Ы�xٕd�w���vn�?K��nc,K~�U��9˸���Ǵy��(�
2�W���:a���ɉD���^��k�?�r��Z��A����>�fi�������f�װ%���@.3���հ�[�)����:�>7LX��!�Wy�h����Ф�����WG�܋�� �g��l���|ܿل�I��|��������%���|�e�9��җ[N&�܂�	馻C�<@S�(^�y5�+2Pe/3ԟ�3�"��B��Sˤ&KȞX�cz\_����N>���p�Q��ɞ\sӮd6��6���-�/S
�4�2A~�v�_����*L��{�pT)%r���c �Է_�x(d�����a�لQ����Ozuub�9w���L����,iz=U	��Ͷ��x�B��08
���Ezs�s�����q=|�/�T�� O@��`t�"�y1����x��iqJ��Go�pz#�|��y8F~�JE�X�j��|�S��x{	���M����R�Q�<�f��9p���NS��J:FڻKKo����궏�D<g�{�ތZh�i�����ܐMZ�[�b�bmI����6��q����!7��k��n�߹��Pr����3-NvswX<�V�������V_�~�g�U�r����-��/W��S�`�M%y��}YnL���-��J��Ř93g�����"��89��B�I|�]\���Ʃ:�C|��D=VǍ�T���D�������7�2�j�$���ظ�$�:m��?z��#�.���~�B�gyު�Hh���=`{>��;�w�}��p..�����������i�������G�Q'٢�t�W�Х��>����Ŝ��ϋM�����'cD�'�SI�W&�]��p�f/��������iEw�a�?|��!�i4̞xkg%�2[p�aC�9f!�i��m��`*}��BQȂ�ݸ����
��~�B�e�YCD%�o����={V��E�2C�QuW�y��s�$������ٛX���G��^K=sȟw��⬝�Vf�Qo}Tc�x���ˏޕ��[�ߥ��%�?��~F&�>O��9I��U�HYVo1�Y�z�_|:���'T饕U߱���ϱ�&��|�v!�(/�G鏦IG��ŉ���u��m���zu\�~�{Ѡ��Q���ǯڍ}HBY	�����Q,�N�#6�G��L����C�<�����k�Rͣ� �ȭ��	9��1�r�i�G� ���-63�5�BBiB��ת�5G��^�"	�c�ܸ�~��C�k��.�^��U4�c�A���f���� v�d�(cw�ۢ��v�V��᠑���4O I����r4���2%&��%|*�?�MqΊ|���y8�G�]_`��K�K꿎��w�@�vN���]�Y��R�����hoa���YV?�T=�K�>/$�/Ù��ɔ��v@	�j�Ps�㙙�W_w~��B5!`o�U�����ʆ[�W��l��'>�3�K�D>N������sD��oUi�L,�����a���Kۿf�p�P(�dW�|S���AV4��ŀ�pV���Z��fO����H��E���J�v?m��^0�M6"�"T��*��6��%�$ �H�?�$���h[��,c�(�i8O%)^���͸�gXE��8�v@UGy-�~�V�y���&7�4�-U�����r$c�=�����?n�\)ɗ�<y�G5�ZI��c��[��0g���n�����r�z�H����(I�5��+F6�����fL�{�6��ȥ3;�&���S|9u�n2�Yy[]�y)I��1�F�O�7�o��O�t�&q���_���T��� �m�5֭�t�f��u��ȳ�?J��b��%9����CՋ�#���F��d�O 7z��~��3l&H�%��L,��̈�{^ȿ��s}KZ����һ㏃�c�e�-��&!}�W�'	�[�}I�u�>ú2i�=S��Y��:,my�=-�V�c�d�&��%�BT^����.���<1~@>�0��7�V�S�[`���vQ���.x0��g"B����#�)��
������T?-�*�?w�ut��L�Q�6ʕ'OԾ��|myjg;�vv^!U�h���nr��x��_���է�V�
�����N�o�d�G�e���O���9IdW�+}�rsT���M��q�
�yY^�Y��n�ˏ�ik�_|�-������JZ�z��×x�{���R�E���\%؉7���0�҄%c
�&�Mby��3];��O���XX��_�k�3��C�_�o��Ng��K�/q��d���yDr�r�P�w�MR�{�+���w�y/ݹ}r�O��js}��[�����eޠ+�vB(���Gx&|V^8�dX�T�P'�E�����M�0�Z�
�U¼uN���� �&w���M�$-�{K�z�[��iiߘ��Sr.����{�p�]؅�[ͽ��%1ߊ�ӱ!|��r:3�T������d{c�1�-yY���6��EQ�L�S�(O��h�]e��P	T��׶��ӛ��*�ʾ.+��#�t���`U�����F��[̯�Y`��5$�����~�E�{�ho~ >9�Rs�P� ��X
k�m�����DSv!��~I&�
	?���eܥ��Q���;���ƥk���VĪ;L���!q�������E�gV"Y�>�>\؝�+A7�m��c�(r���N���
7��!���%\.�<(�R����r �A,�*��C<�ϣf2䈙�,gf���r�[�IJ:HnT)Ʌ{��E�D �Ő��27>"X�j�6yYN�y!�@W��Ȗ����#ܕ$�(}�6O��e^�rԞ�z��^�D�c4�:L�t��� \�l]5n5�>E�o�iB�p7^��&��&�u�êby��ѓt�� �ͣW��# �����ȷmM�+jI�Q�(C�>+�lgf���u�f��(*KsR�_^yA}j��;��}}k��u����$jB'r̔�g��|[A�J�9�6�?�؍��*b�.���1���$��$<����2�i�ՒS�d���rN\�Nugi��'[���wށk�S��tzu{ �m���/�k��>�d�\��^��!=�൵�`��'���d��Z]Y�_�Ժ�[o��}5�S��#�)����H��`��8`c*4b��|����1�}{��].��Z���#��퐪��)1��z�?Vױf�K�|D`�K9�V:6��Df��o���}�b��6��5S�ȅ�~�s�Wb�$���q�¨�BSS�����W\����X�;��[��wX�Ωuo���8�a�¬G�;�A����d�v]2��9Ju�)�~�A?�b��S�6+�RqH�5���
��Q�>�
|6Z�Å��
�z���	òq�>"�w��0�p����:O�Q�R�/�ll�nG1\q�c{6�U�&��1���V�%{�q�L��y�5*��&�G��y�,��Z�M���C¾,C����~#�`m�[�C��߃c�[�V��i|k�m���y:�j��v7�i����gI^Je�(	n&,)X6����<�o��Fy�;�$�NNO��΍r>rt5ͩ%�V�T�|��=�4��d���C�{�O�����0�]��O���Aa���8�_���H�Kl������ֆC�_��R"�R\��p@���3=���N���I$S�s'�.����2�/ ����L_�>�1
(6�w�;TH؝�=6}��<'�Ē��rT mj˾F�:��[a�)k�3j_XVM2{ؔ���-{^Ha�LL{�fΖ�Ő ��U##���ѝcr�O�p)��g#�<�=�"d�������{�?�ǹ$^ύ�l��~E�G�����mm�����?#킛�AFePH8r�f�f�-wG��[xM1�̅�x����<!�d�;��%����v�H��麪�	.����C�bD�L�ԧ֋k��b���5g�2;{w�A�
ۚ9yy�&&&'�kk��i���}��P'߼�w馟�O�z}Np}��i {�����AZS����|�SW%�h��x�˗��<����{6:���nsb�5�JvT��Ųq+[a���$�L<��'
�V��W_	mI�oZ���d�\���^�9p�����#��?�I����u�2T�Q}*�!aU���y��������G���/�w�F���a�U���[��_<��6���u�m^>������ޜ�|)�>��Ҥ��Ȍ���_�g1<]K�)�A�����}�Bdy2�GYYY�a�Q
x���������ce��gB���K�����=b	�).��5�z���(�2V3-���s��\���P����ڿuv�k�h��M����q�-)���8��!��a�O� ���ͪ58 m�� ɶ�u=p�4��vnu���~�G|�"�<�?�T@�'!��݈��5SE�S�2�&��K�����Oe��H��/Ï���캹�z�/Z"�4�_����L2NEE�������G~��{o����k�-4ב�a�-,���j�T/�0X�D+�W��O6�=x��[Yt-�
JH�2/5!��٘i��sޖ�aV�`b��O�����K!��d hn��ş�
��%�%�V8D���;��F|N���p����Uc��_�Fy��9	v]5@������m�w���#�N�u�*I?�SܷY�$+H��Þ7(>te:d@�;��x��A��M⼐�T�'�j�r�0�E�.#i�΂���O��)��F��xٞ#�~�N�H�_m�${R%h����^��=���g j�a�a�4�؅��bHc��{�ۧ�f��ك&��� �χFF�ǌi�nc��"��Ӂo&+_�����Ud�G�Pg�c�dg^X��9d0�Z�=Kkg�;�߻|A��Ҩp����'G��@���w��RU�lWU �Aȳ�S���`�;,�X��[7�m4��'���w7=�/
�7iP��5�R1��-O�V����w"Ք��S�nM�?S�K=�?�!-T�*�#�\�S=�wf���^F�9]���|T���k!|Oy�f�����[�暽p�N���[:�\��%3��i�8��$�-)^Jp1)�N��C�����y�=�b� ��6HY(C�z辶�5��}Ն���p��7��0V뎹GN���xn�D��3�^H�٦�m���f��z���.Ei6�}���'"�
AYO��W�p��Ԫ+���������v��K7Kn��*���_�£ׯ�'�L�5��gv���Y�$����P��P���Y}���w�z>�7	�Zm�Ql�n��D������@��m��yQ1$)r�	��iS�m���9� do�f�5��/V����chȊ��w�Ą8��}.����@�������6����-�4�)�eh8�� ����}�'.q|��]em�Y�T��k�5�'-�ؕ=Hf�ȕ�3j�R��_�/g�딾�J6��#I�}�@��d����p�y�K�wq}������j�g1��k����A$b��$��0D��ȈVye�|O�e, ��6ާT(�7�L���������2$2�����W�? �8*n�
}�u�@�%���'��b�����H�j��G<�
�J�������o�D���r��1�z	��x��,�(+ߐ��;�`{����t���a�s����g1�c�+7��;w��WH����ݮ�A���A��𮡜�h�[0��		x>�5�f��v�K�D���~�g���d kw�o�
�Y��wܬ���m�}Z�)���+-�X۴i�>��G�z�/'5$��E�v{>m�[r��j8�*6ۓ�M>z),pteZSgw�z��˵�%O�{� p�R���į4ֶn��d�'�v��������I��dݛBYP���-9t+�K��~X>dV �6� �1������Eڐ��Q�/�/��hia���EuFs�6�ttt\/(��@�5�/~�E�sA�d%�B�^j`pp���6�P�����Az�래a�> l�V��	�um���/�k�>u/_�UK��YL�	���H�m�5^�Q��7��q����K�S�$�ϝ-H��M������N�ǙE�k�7"�u����ȕ뎓����J�
\�9�x�E0s�5���UQV�m���ꕳ�Gm�#(
�-I��A��o��eݬT��a<z��1����%o���p��sh�w ���6t�{FF��G����$��i����w�ES[�5�{�b�:��;E
��V�����-�J��G���y�`�I^,i*� �� 2���3T\��Dy����OX>���eH���A����[J�`="`:s��)��q+��r��,���Q�W���i|P8�0՝;�#l����-.�N�u\���'��ld	4����եߋ�s+h��x�ro"b�}�e���@������Z�Nc"oJ���A�7��_�����0���[���1���_L!/��Y�MGH�	��䛳� ��Q"��vdo�{�h����$u�Q�@.|_x%��W�q�{w�qN�I~�hM�1����O���d2�r����C����A��M���Jb[41~:F�T���R�i$�Td�����=(�`)��{�
��G����\�]T�:@�����r��^����aPY�LͲ�c�އ�����<�}<<t*xQC����#�!���r<:\Rc��;W,*����X?X�x���<�Pc%.�r�]�F�;^�.�Ǒx��b=}77]�U�y���
n������'�Ӱ�wx�R'؟؋�h���vc�f��Q<����	!fn4`c5̑�$��ʳ��id�$Wɖz��^m]�p(w�GX�\\@�1��b��k�7��MuB�hZ��_qcأ����e��>Qm�DiL�������f��L���=UL �N|�4RgV�������`�8���Ʈ�K+��/y_��7޷{�A՚�����e�:'Eg�ϑ)��"��S��>�tYt`x�"0j�!?-�����V����@�HǄ��x�s�S�ٽH�����4�#2��m��:��j$�J��L��L�oݽ�����"�v��� O+�Դ��My�ɦ���|\�v���q��b�x"��FtW���nA<�7�4��^��]�N�ߨ�(�Ҵ�I��������wn�̧6i�i�pu�.��M�V��I`P�08��H��>�(2+|>��=���;��7��n���N��8[��,�:��ੲ�M����2�6W�g�X�j� ܬ�C���Z�b�s�ъ!��g{ko�����";$r�?�f ~��\�6�u*�JSSS�ƞqbr�İŧ �j�<=BT��U�thb��N���ņN�#�����GL
?ˋ����t�W=/�:n���Ȫ B(7����7���a_�W��&�06�c�p,Ҫ�Za���v��oF}���
�Lqw���)�:2�QZ��9:6�_[[{�`L�~1�,�K?�tw��&AymdB�cfd��R�S���pݦgN�?�x7��P�~�Ɓ+d?�ɥf�|ڂU�}1����SY����5���턦�������W��f�F�jFx����!����tL�G��W�*�PavB�Ѿ�{�U�g��d�(���Svf��n*����뽫ч���F�-O�ǆ! KtKt�n��/M�/�~կ\��#�<����y9��n�f�~��M_�P�η��~oL\ϸ�߫?ݪ�f��v������%��	�d#��I�ɛ��1!MV6�>�Iyԙ�8n蔼�VdV��
$^5��G��������n:!jp������+�r���'��I|����RK�O)�2��>[�4ҼE/���)W�/���}���2�L��
¢
x����]O��8�Pm��Ɏ�\�J��P�8R��S��bp��Kx�^�=^S���6���?j2[�D��Y�eˑ����Q%��_�����g�'��y@)1������6
��xT�x��ݱ~�D/�	��KjW�Rzܻ$��J���j���(�yg$c�n;��Bf��'��1���s�ͦe-��T���8׽�S��������H�gc���5��I_S	a�K<���e(���T�"�{�=?8?�k��G�Ee��,�rI
f�lm��Q�d�;��~���+F���ƪ�Z5|]�N+.��2\A��e|K;�K� w�r.���C��<�a?~SHI�W�Sp}$�J/����p.u�,C�fW*Z;i�(�{���p��ȳ�-K�&��� .��)[>==�FH�u�h%"c��$����y����-yړ�-�@[�k���=�oiy��sf������y�-�z�=:~��:㱧\,JN��;�/�WQQ�sz��CЦ���`��3����{����#Ň>L�{�f<y���_q�����3�x)O��[<I@�D}�z_�4��w����;���[H}�U�.�ۼP�}5e��wjX��&�1#+,DG���ڄK�d��2�ζx�1L��%]����������q����z~�a�R�1;���}��ϩh�Df?}n�����Q':�v��R��)"��p.�q1i�	ͩ��b�J���&N���D	�M![�����~���L�t���a\pZ�h������{���D���!x"�+Ap�(�pY�<�e���<y�dd����9�	�l7���=4U�e@h����#��w��DSs���df^qژE;��YY}��r���u_IL���a�g}q�E���#R%������}8�F�g��|�W����4�ЁbU^̜azf��X��苷Dw���OE�ʏPG�����#�'�v���O�����e�v�2w�����G�ҫ�t����Y�Tf�:MY(uq�<jr�tG��$΂�}��he���f�\��v.�+eK��Ǎ��Tu�G�Q�Oyq�fIC�(�L��x�o,���)��x RA�ٷ���RU��$�^�Hr� pD,���}�%�[�(0w�+p��,f��3^pӪm��E��^M����J]���ݏ�w�Z�ͫo���)C�ٵ
0u�����]�4���~>��A><<<Vb��p�Ly˄��|�t8 ��ՑlG�Rin0������)%�uB-(���ב���#���t��Ru�|���+L�1;��h�ӪaCRg����뫴^����wno2�P�V���MI��k���8�q�"�N��u��sb��bp�}4������yv�}L�$�[��'��O5o.��z��R���65RhYӒѮ|���~2"�o�\h�_>P�_���i[���2�p�\��@��b "�MJ�� ��jU��s��P	�(Y�ʏ�M�)��)���]{1����ڹ��J.M;�7o�c_�X�`_'����Pޛ�&�u񥮎*==ݟ��R�hz}�m@Q0EUWW����/P3�s�p\^��Y[�Y��A��Q
2&H��� (T-�)+9ާ�TB�����SQ��j��~33�G�������1�,����;l��ᛓ�ׇB�~�Ҩ�͗�+�WP��y/��v����Y#�5�.���Ol��Ll�ҡ;B�,2G��܆C�%�0��f���6������S�	/�;CY89Sm���>+�T���'q]R'r�R�$�o�}��[",�s��� }�����U��;���w^�E,p��HuHF�ܲ��+ϸ赁�F�ߢ����<pJ���m�83)��l�9C�]��Y�L�@[I`R�w�uk'��pe��z�E�ϭ��Qb�~+[z_9�癭�?������>���"!�"H��J���-!�ҍHwKH�t��đ.��Н����{���ُ�zԳb�9�kͽ��ח�!����V����&��}�v8T��Rr[/ϴ��f �������]>k�mAro�@Y��IO�f|�L��x�c����s��\��č����Ɲޙ������
��L�oW�{'���2an��ܝ^��XQ����@��ի�I�0=�$hu|qe��
GFN����>��Ņ;;;[�T�=>s�H���7w���P93yId�AB.��9&�_G(�3P�!!X�dX_�*��|s8T���W�N6$<��L��������4�@��N�=NW~�𹽿�Ә��X{#���'�����͟d%��~��	[���R)2/�P֎�Uib��ob
9z�Aٹ���\k���;9���8���׍Π�����n�`���&=���O!��v.�U^ẫm�!v�w�Ls�q��,l����FM�1�w ���@Q2yab5�oo�iݔMRI�r�}�3��'�f%�U�'&N���u- C���3���<�XJ�ڵr��;1����굧�Ѕ�>t}�������퇯#K��P��@�F��Kh�dߥ0���fs��Oɥ#�5*�f%�L�Ϙ&�|�����y��_�F�#��݀������e._H4�Qt���
~~�N�v���?��#��%�w���g�%$)u��3%.Җ���@�>�2�@��ǀdIBBB)e�{��~��e�-�-%-�ee�J�&�%5ޒQ�&R�>0�����ru��_\^�Dw8���h́��>��\�z��U�"�oL�ޘ(����s��&"m�F�v�/LZa/輏"L��ƆzB���11�
�O�ϥޢ�ƚ8y��H�|u�r8d�Z{F�������ؼg���'�S�[�J���m�ɷi:�<z����wJ�@̱���$�v�����u0g�wg�(���d�Eȋ�(CF|�<��Ȝ#pK�.�?�[������(뭟��Ò�b;��I��8�4��YC`� �F��� y�椻or<�LyĶ������X�H<A9�B,	�b��of��߽ٮ����{�E�d�[���վ�����s�׷{�>� E�Nm5ʞ�b����X�`��U=2��J��o�gd_~��}T�k�B�y	�H��R��Q/jy�Szv�G�_�P��"l��cض���/�{#@�e�E
� �{�>M��[��v�`<# 䖺����[l�@s����he}����P�f�7QCwߟr=8މ�{�p�S���;����+�Y�o���F8"������F}w��3��(�I����H��S���MR�-�,Y�P�h<}�ڮ3����8��}>�s��xG���Pkzz쌡Ȉ�����|�t���������n�CE_D|�ˠ��0�HE�u����$�>z2RJ4��bX���jd[����ǝ{�=wC'�����JlP���AZ}W�����E�i�ǔ�B��ժ��� 5�J�6i̓�b�,w�W��.k�><�U�pj���7�B<R�ጿ) DMMMw�����Hd@ɗ�`[�P�[|bo���g��F�?� ��`�������FZPwD�}��m�pm��WzǄ����DPP�߻w-�����1���>�
���Ύ�q�5x��֣��D����"ы�i������p'��s�a��#��,~�P���f������)�%H�5)���ޮ�ܨ˜\UE�H��>j�޺��>>M7���rX/j�d��e��7�x=.�V߆��J�7O�A"�޶����tqqQj'�4�� <�2)����Ν;l���,�&��x��tyKC��0������]�?\�8̌��r>F4�Ӭ-�H�Y>Ackkk���5x$�j`]�X�M{b0|""Q��`@)����00R�����ݿu�Z�/T�b�aaZ��W�y������Y�=W�[0�v�lSz�_�ZL�].F���1j��0H'��::���T�����d��������Z%/�?�\���e�৑�U��U���9���B�f9��}K��?Q���c>��z�����p����7��@�Q*۸��(��������B����A-=}}�@s�@�P]=��X��oy���9S:�1�ߢ�ˀ�l1���Xd����x " �/}: 聓����B|G''�хg�dd��Id>c��]�����j�L����k��.�iK܄Y�Ӡ�ِQ)��o�����m!w��wD��rpPj��f��P$�3R߽	xRz��H1k4�ߠ.�h>!�'��P�e���:�]��M��5�;�o������.�A)�^	C�6�����<ߔ��W�iyG��=�=S4�3เ�n�ˑ��G�0���XqG�VF��R6,��G�.��X��0;����Բ���i���f��7`�u�M˜������[��)�g��xcĴ��`�A�o{j++	&��7�}i7y���(�q��$N�!�RPP�n��D]D �ϽD���"51����C�bbbr����f;�ԯ���*V��.�	�����X��������r25��;hfL���v1����i,����Y9��8�O���0Hw��_�� ''װ��8�������f���"`����t*%wy�z�6֪�g
[H�66,�yn�0��a�^�i�FA��|tt4�i/b��>��|��w
��jA��,��>����)����1!ǃ؋�����|�*(���}�ؼ~�ĕ�K�ϳM��^�Ǒ��0qOL�O�w'���&����w?� D�T���%9��-�F��G >����߃��0_�b���� �gb�c��.�7H�1`500x-.�����+k�xu��U����{����ρ5���'����Q
?�咈�J�NG�ﱿ@�~Y��@WqYb*=a"~sũ�Yy��w�:� ���&�8@������c�7c9�T �ѽ�{(*'��<�Rw�g!'����uy�(���ej��^l�������5gG+��$����^B	��s��)����\-��e,�������Q��uH�����@�c:��`aQ�!�|<���>���e�s��)�T��Jnl���h���񝬬����yZ�9 !�YY�>p����������@��@�zUK�p_^^�ַ4eUiф�j���/>L�����7��c~�yI͢���?0%� _�8j��z������`���;H�\���DX=b�X	;>���<���; �f~�&ce8?�Z|�Xcy�e������>y�Qq0�o9b������l�d����V��QdH21�`Ee + �h@�� ��IZw_8:u��<_R�4a��M��Ұ��m2R����uQgA�z�&�ņc- n����W��Џ��U��{r�e��S�c�!��X=�k�Oo����|ҶQ��/��*u����ycu��(j.����B�����AxC���1y	Ւ���M>����_G���i&0<�����C#���Nŗ3�=^e�Tj���tݍ���b���$2������x��
�<��
2-�*���lox��z�(5'5D�V(��V��֗��EG�W1����m��Дs&H�Y6��)]��G)��g�?�J�'������6v�!h$�̼</06�u��	v�H�\݆���"CM�|�Y}�.C͟*�k�2M�Z(4��4/0PO�W���
ƎQ?6��<`PdT��A�4�>U/�����:,���v��1��7s�=���~(&��활*,,��#��M��_.%T��R���Cו�"wk���p�~�@s
�l�H��� �W��m3eu�.���)!�F�N�ޱʑO�=Z�4�[R>�X�_��5��tDZ9��,����ga;�� ӗ�}�9;'N�K4?����OǇ& ��1BĞ�t��xzz������r�h�.T,$:113��u�~+	~a]�+�6\W�τ��?���.��~@ $���ڍ�Sd��J�,Y&r�Rڰn���ŵ`#�'%����������(5	�J�^�F�Je&k��cn��ǈry!ɫWB��ˆ^�%qv/�{��A�&d���Q0�8��= t��Nw��(�mm��)X�;FE�YyjY�K�/�)K ,%�I�>(ۇ�Q��de=��U�S8Y�?�U�S�:^�?������W-p����z���>c��Qxz0�.w��^�4vU&����H��	�����{=`&��ʣ""�KKq�ѕc�y4j���	�(1�Hf��vO7�~��َ9��*UZ�=�}p��`ra���������]�i�_1F��i �-m�I�</YY?766�"#9e���7,Y��<���P��38��(&�����P���M��M���6�k��s��}@������%�eC��αo��Y1g�������:�
:��
�n�F�j,Q������ E���$Q2��azs_J^��B)o0w��b��}W"�����Ì��*Ԏ����W�z��	
��h�#-�9.�>��م���l�q
m*c�+y` �a�<����V$| �`}��MF.3��`(�7`�n�bs����.Ƕ���� ��Om)���z��Y�K�&���4�O.��txr��eP�t�1@�6f�')!��(� p!��B�Pʷ��)|?FLq�^�������bl�a�U�6ݟzQ���xӉNk�St�/A�	?ොq�g�?�5������k���G���5 h�a(�izF>�>g���>8��?0P8&!�  !!a�ؘsC���_�D�����Ȱ\�R`���	����-���U�V�(j
��|c1��9��m��{a<85g�ݷ���OL�+_���N�[7 ى~eN��C1���н�?`p����G���p��M�H=�¦U͛��E��~��C���� �e������5K�X>�U��C:�G� / 5b�ajJk�U��2EEE}��b�͢�=��ꠊ�J P@ ���qC��!��Q����b���n��p(s��bN��멙l�WD�(=rt��Y�^��V�]��s��w=�/��� 芑�?����IW�h�_��	&��}���{�S`����Ot�⺇.�tѻ,�w^V��EY��<�;F�L ����#���;�;��֏C�t�sz.��YY-�8{Р5��nw���k�Aƥ*5۝���sQ7`����7��K�o�Q\A�2�
�~���{��-1B���F|Y���S;��~�C�_?J�yt�Hq
j�S<5س�&��_����{���Ǌ�O����ȅ�JJ�g>�����Jr�
��V�Y�S �AG�y�ݽ	�w�N��'T��f��cu��$��Ey�+/,� ����OK����(Pݕ�+o��d9�DTD���uS>����I{�Iz"��H�&�TҒY(���d8�*�\�"yjNz��-"\�sk�9��E8:�O��E�`�s|���ԅ	V�NY����,�m��?cK�`�QX�ڒUu-�Iܿ(w
`���}3�g6�^��}��U�	��h�^L{1�xף%�7^�yV~\�iD~���6$|�fT�����J���}�[�y�5�� ��O�f�-�%a�wv%T�Bf�_U�I�j���Ė���a�����
A���~XU7k7����ZW���� @W�#�x� ^�S�`	�z�>))�(Hk����ӧ�� ����L�핿/TB!���0��H�L4d6��	��i �V5��<�Zq@�%G3����xϰ�r��9x\f6��ȕ��W�ߣ4n-aU�r��+�}��q3ff�o��n���j7�����4f;j
&՝������o�O��UU~���A�E��c��˿�/+9�i��'�#����ӗ. ȗF��O�+)��_�V(���=��-/O��E�y����UT�Ć#Z�?���~`#� ����(x5�F3?�xBvp��@� 8�x�xV�� �#*@0!���d
Y�P���*�<�SU��4�̗�D�hR�U��W���v������g,��;�K�#Z�d��s�Y���^:r�{O���^�/Ŭ��9U�HX=y-�}�q�Ipt��m��u��rJ�K�xq©B�ʐ�/�:�r[��f,;���TtYvJ���	D���f�ܮ#���΢���-s��F��no�b��b�y�ʺ8y�����g5�b����jdb޵Ї-ɕ,��=��ő�4�e���Ԝc����/\�NM�׎�~�Xw���?N�Ǌ��e����@j�t�Ç9��"�A-i��Ɔ�D�#C��:��ĖٞHz��u�����ݜ��b$��F^?#|Ѩ��Ja%����)��#���uU*�YŹ�<� ��@Ǖ]Y^�	jyG��iϤ#�[��=�kB�gaGs�z�2������������ǯC����pͳ"����˓ob���k�p�� ���')�_��������\8c�Zh��p�;i�@.� �����V��`�&�k��1�8hw��ƥg���n�ӆ�1�n�;�y�϶:���� ̭J�c��_C��@pyκ�_k�U�(bp�t|r��F��f�6///5p��9�׭���X�뵷��I�ۉ����W�Wh|�b9n6?���p̪;E�����}�/{��UޢK�L&��&r/�I��B�tw1�r�Z�u��>��T�ecc�@�_��˪�R��c67/p�
K�,+��U��(�⡅�|� <=�<�u�I����S�_�M���D�"W5]^�
k��Q0���i4������>�劙my��9+�r���	�:N{=,�'�4m�$�{Z2�Y<&}���X�������cƋ��ݳ�n����0?�|<y^ɨ� ���mbbB�E<�G�X�+�=>��6:x/mAMʐ��i?y)?Y2�I=r�I.e�B���lIN��Ą 0�ʥ��/�^@�߾���-�pn����t
��;E�_W9��@4��71�IK'/�ep�?h���cq.JS�9������.*Þ�#�d���V\���6d.���si��ۆa�R����c���jf����-��"��#PPQID�ie�A�S�lU��W�D}�����i<���kg�/ق��(��/�*�=s��ڮ�������B�"s���z�M��/:��ggS���m	Z��=]�|5����J�Er��2���>�u�S���ٍ¹H�����7+�\Ը-�B����j����˖rr���a�,.vK����� ��=?���, �z)+#qF��-6�2� ��8��-��>W^e]�=��h�b��w]�,�w�-}�8V�q������v+*
���>I�<��X+��������d_X��L��6�hf
G9�����ŉH2>W�E�w�\�sC���
وI-�� b�+ ���"x*+��9jftMT�Va���4>���tc�g�kW�V>��
��ֲF���C�(d<�a:jd` ńOl)fk[���)����D�=�/^(���vq�ǃ�x�+���}A^���ҥ�ei
;E��"�|K*�)��˻^�����R�zjQ�baa����,���o�܅i�����]\N��41�}�&0���Zɯ&n�t�^8��Ө������u�!H��cV��5["�ey�����о��?>�}e����w��T�/��'�C��-�rG���O�Zf�ΎVl �c�<:^$�w�X%7�l���y�k`�R���]O��1RZ5�J.�(QaRTTF{�H̳�����څ���^�ac���ngʑ�A�P%zib���qP���ά�Ĥ�~�%��R�N��?0���=�>ZLeF��@$IaR\\ �2f����	�Ň��AC�M�P�5�k��ui�iFԵ�����.����٧1JfI�Ne��3�*��J��s���~��ھ��VDY������O�H����Y9`����u%_���UTLg�{>#*��"�o\^L�t:1)�`$ @
���:9qI�� ��1����H�Pk�aSJ|U276�[)��_]5��헥������e(���ة����x���E+]@W����VT��0��E�3 Q7 ����1(n�o��QVj��/G�=@�&���}�/l�����6�Om�T[�țZ�W,� |
D/��7�J�k6��X�_� Hs�{�YF�%�o�����W�f��)8����r�^�� a�T��4ŕ�
¡�6�G���
W�Uۀ�D"�x�9+�,��)|�nUc���?,���4X�eU��䝜�
4�8�k����|����#xv����%0b_��І��y�j"����4
�L���RVV�xv���ӷ�$7�i{���
�N؈w�4Љ^�E_F�����e���m�Ћ6Z��7�F
rs�=1y��Փ��!�`A�����r��hFr_���nU퓘���{^�Vwl�0֔���426&�@��)y�3퇚2��vL>\��d��bBbs:,*Pƽ��������V���7�ǖ�B���E3������R=ǥ��_�ж~����!��m�Z�Ҳ2#--�_g������ �:3
�
�N�Ow5�Kњ�YY}��GfUK�\�G'�q������݌5Q�%?Yj�NC�@���*�񔍌����"�e�,��T��2�8D�K���w�ხv��㸼�f���=@d������:f��G���d�%X�22qwNA�v^A�$dwCì��u4I�K���[o��hH�ք���§`�\(���t�A�ոu�(B�)���XN���4���`b���Cȏ���G��H8mŠ���S�ת���N%Sh�ԯ���~�ӣ�޼��ap�I=�&sA�"���ĵ�CG�,��u�z2��)<�PV�]��IWU0�n�tS=�1���&m�.�E���U��������
��D3��t��HS
]��"�M���2=t�2�a�_���/����f�ꉳK�7[ld���;�ϖ��V_���5iv��Ә��x\��]NW4�c�$J�G4�^N��nl9�
@n�� �oĹ�5u�3�e:�U���=��k��w�B�2[���UnT��UpL�[���6��,�H署o檽��3N�ܠv��$���b�
��"т�9E�Gi�f�:��x��,$+�F�mk�Ҿ��WB=%�s����(x����[Ps������F�.3W���u������A͛i`�-S��4v���ȯ�V�ꡕh�"ٵ��F59�����]Xz�=W���VT�z�qxT�$�> ���^��7�v�\�bgU/��I�p?=�"��ʛ_r��n>8�$`�l����ez��O����?�&AH�7���0��vg��k(�j((G�U
H��+>bA �VP �9�}����f������u#I<�	��g@gdt�gH�ONO�;i"�M�B44�E�*��q�[YXH����f �<?*8_���0~���-@>
g�)R=��:���}(���	 -k��'b(W�P��WӨ3�ݘ��*bO�O�]�J���U3~�@åm>�����i)��.x$}մ79�x,��b�|G\m~���=D��y��UW ��1�����3̑���(���S�L�����
�R��QK�p���G%.:�5��	������B[��̤*�w���[��u<?��1�Vc��1��';�K�4B��YLYÑ��7���p�Fr,�]�	���[+��*0��ԫ��頼BH�z�쨪+pS�)���O��Jz�s!̓}He@�TTUA��޷��b�8/��w���p�MN )7��(���b��xu���zg�:��[�]��b;��E�#����遡�����m:Z���xǌ;Wj�T�s�g_�"!Y�����	�p[�Nގ��e�<�Z���kk���\ ��њ,�H`i��E;+��*...MƍZ��sl2n�'��~}?[G�;�G�Ri�?ފ;�*0s���������<%��,W��4�Y�Z�-x<�ŵl� �UmwrF����2ט�{���y�20PH3YJ��d��)9��7�B""�>�W�,à�>�?-4�+��d���W�>��x�.��u�W�Ѳɮ`��fc��4j�����%�4�;����N���(��Fff
\��&h�&����*@~�T���h'�%����o�bl�2dݩB�y?���͚Jd������&�8��s���^eR��j~��Ū�*V�Ek4��2��٣�`����,PV1. (��k���R�����Fp��ڿ.3�$Au�]�iK�<���w�<,A��U���Q��"����_�����5@R�p�3A��z�a.B�x�ݹ:'G�x}�a��mzͺ�F�ko����Q���M?��@�%����N���d a�j'�pIL�w��B�H=a�X5i�'}��`L��w�h����5�t=6�z��{��B��+1aS��
2������ō�n�~���|ౖ��F�A��]��{1)�}�+y��55jyyy h�V@���{�����WPw��a�Ǻ�g�������v�,�	8�
I�ɊYh�v�{��~�8�\�
��$�PS�Q����{�@��W�޾y�������5"2�2���xu�����(p[�� *u>�|ՖHiT#ΙcC�FE8H�a�����d2fj)N��ܸ���V�;S����%%_��X�A���:�]S��@3ն�����0�ɓ����C�5Pj���ސ���w�sܣ֥���-�_]7M^��z�3�R���ۙ3�-��]�ܪ�A-��L6���מl���+� W��ӫ:��#��><�@�"�����w�eM�fLh��5�� 4�/	5�]����$�W���d!_889}����奤�@ǣE�=;^ǜĸ�9Rj�_��:�?�9	ss�h;�Zb��]�}[����G���������i�{C*P�����2�MK0-���Gg���ʦG�}Y	�0���[�j��ϔw�T��0i�S]̤��(� ����m��b�5?/`�M��98�'�-��3w4��G��, s�mK;;�<Woӕ	��7y"��Gם.G����ʒu��PZ�%�(�7�fD:ChK�0�����������Q�nګ!����߿���Y2���剛ן�m &&4Hح�E����#�*d�qQ��f�Sv�@2f���RN���A:��Z��˩xy5��.�M��XQ\6��P��Oh���{�����q��+�s���v�v�J�͠{���q�"��J0� $����9::����i��fP���D���dZ���Z���z��#�ZE���U��+d{���b-�r�0�C�1����r�>K�{�P/Z��Z��� �N�L[
���+��ؙ��j܄�1bz}yy�W�nw"�:o���o�#_�*a�<mM,v��@*�@���[�gK�K��T�`7�Rj!ϖ̯���Ԓ��e�����ި���L3=}�a�#�t��Q�Rg����5�U{����MH-�ġ�okEn���&X�%�e!�������ْ�ВF�2�Qt�Q�	�"D��)��hB^�t�3ri>�G0�dXx���>/E��[��/���!�#bI����**�+��\�D5e��d����،��b��I�Y��2�kU+`-�rO��W:9����k3���Y_�u�zWY�XW�SD��;�{�x2%����V^q�r�7��#�(pqp2�r�q���J��,���-@����AsQ��-�fލݽ�,���os=�"��H�ϰoEv����xS:�ϴu���N��Z�#�s�	]��OQڀ���"Q�-�c�I�ÓӺ0w����o@
-$:�/����g@�����]��?�����T�}[�[b���ʶXy���F`Y1K*f2O�E?{���?%�g�BXׂ���%���h������v��q�r�>�TC�W����z���Ԁ���JM�:0s�d��f�n`�s�ׄT�d�LLֆQ��1,��h0���ɕ��N�����8�� ��7Z8��͑IC�n4d�����ȗd	:�|�C7�,q�g�Tp8e����"  @CC���]�g�.cl�H�$��p1�<�m�Ɋo��W��Y;���P&m�[��><���.��:#E�U#^��H�k��-�'� ��b��VO�Ji�Ւ/-��r��l�:l8���f��iV�o!*þL{\\���-(�.����a����Q��ꥆ��%�=L74� ��q$��
~�t�y��蹜蟂�1�9�����T�SU?�W4k��%"4?�4O�.0�+3��c����~���i��&�l��i�P^.~G���!��~0��Dfo�7�'WUqd�^%�׿7�E���
���A�g��֣*A�%����h:��^�Z��0J�uI�!j̬<\�Ack�U˚�et��z蓌1b�EP S<��z(��X:���r"h��ړG���r�����j�V�wxH���[���xw�v���D����V| R<�`K�4��^^\�� \5i'��-�׽��3��vE��t�d���dε
>I���+<N���k�Y4����VH�E�O�c�!����Zr�{��RM��h]vvv��"���D��+(D�h�}t��ԣ��� ��hn�����Փ\]���sJCMF{R�KWƣ�vFp/8>T{\ٻ�<h˜o���%P��:z͚x�%�r��=�v�N����H6?�a ����4e~:T�? [}j��pّb�����}�O����e�*���n��7��?y{��hX���i[�YmYʕ�*�2-�''!x�z����vo�֞�sqY�$I�$�?���YZL�RTi��׏��~̤�qB�����n�����$Y���uԋ�m�F㎖��{�*��ü�	L��*�?+� 77w�w"],����,@�g:^M��R�������|0W�F��t���Y��*�%#��#."St�ۃ������:S��K���\8�����5�������k��67<g��pm:�rǓ��Z8::��o�X�h �h��T��T���ռP���c�ex�}_������H�����wnh]]��� -���P%DOO_d�*��BD��X�� P`>�|��� �=��B���wFaZ��n����_�Z#S��J�_��ț��5������{���خ��f�^^^4tt��=iO���3:���D	�j

�fgiU�zu�4j��2* �8~t��"A��L��Zہ�����~�l��K\�V( ��i�b�}��c���`Fȅ��R��q��G��v�f��og�/B�Y�Ӿ�w���\e��F���`V���Ȓ����s�[\J�im��b�(���礥�SPP���������@7� ui:J��/egW��f]ee�ȏ3f�`��n�������Y[Q�ӝ"-� Vm���`r��<�˥u�PhvN�M�퇙YY��l:��bҗ,�a�?�DU��L�ǟ	�T~� �5O�T��n� �)��:�w=��٭`����֥�-b�l�|�}��)quyaa_++���U,h|�o_�v ��&��40<|���/��)sh�z�����E�?M���Cj7G�Q��ja[��ܙ�^ǏH����ŝ�p{��tS�hqq����?0ǝ�@���e#a��%6�|u1˫$�n���k+B������DO���q}��x�uK�4��6"�ێ�Pו�c�>~�<>� �?ߙ ���ܿ�	�ד��5kS�J���rҢ�������Y�^���;�E�2�'���֭����Q�q5���/�v�`wy��ĄX#���/���2�����2�V)Ě���/����¤�:_��#^�7Ş�6+����:�g���ǆ5_��z��"HX�i�|O�����n\�_Y�}��g�f^�-��B1�7���v�%��H7��|r�yLY����&_7��l��}v�*,���#K{�WZZjğJ�s% e��ֳ�d��w�7�����7��YlO�e��X"��E�䭭.�eg����	X>��n�Ꞅ�ǧ���~�ғ922��ݞ�g~��ʐz�?��Y�#CI�X��1��������p��&���׀>{_m"Q����^�-(f��	L+�v�7�J�}!ȼFFF���+��]����	������4?WII��y�3�rw�Y�ةli��LDO/鼿e��""��z��ٞ���r���� FB�$��n{6>�=t�r��ü����L�8ρ���Cۋ�	g-
m�r�Ȃ��$ ݄C�.�{q~��@�4:�a�DbX�,������C�	���IÅ:>f5��>�פ���a{�^t��r$�	�7�o��E��	�.˯�����p9��>��,X���$|W!_-�hT��oSi-���˿s
���3�烼F�+�b�˫�j!�>�-�HY�WU&?~�|��Z.�Kc�,��>��pXH��������24�F��X�RI�sI<�U��Ŝ��B}�:�����\{��j1p�W��4(���&����uj��͔�� 5����Y�E�&�4{:�pҹ^�Eȥ�)(�OY�_��Ž45�����o�r��B�v��a������!�u��1[M���:����?�q�=�Ӭ���uc)�##"��!�� ��A2'� �~��rJJ���xtJ�ޙ���0O�=j��%���f%)x'!�u�U礁R��j��Gm�(�(f��5�4+a9�o!�CM�B�����{�G�(��k�����9 R%M޿O��w1����[[[%�K2��Ur��nt@@V�D-{���ή�r�q7S�� �[F��ƻ�1j�Fook���LJK�l��Y8(^�-�������d��fN�ن��YT����"vA���q�n��v�/��q���cP��\HI!s9,#*�QMmX9�յ�L-�6Z�{���,����'@��տ���)GR41�)(�[��ܑ&�ֹA8 �I����`����e3e]���R��v'*Ǥ��$����R�
m�;���```@�P����/���%��t�õ�J�B������C�
mN�R?��q(��G�pyih�8P�_ժ��S.d���8-y	va=jC�cBӄ�S e�����S�А7�;p��&" ۃ����w�p:W����3���I���8�c��hH�������Ud��w4�o
��v������yA^�}�Uo��>8:9A���/��	c[�ݟ�%	�j%��z@^qs��*���Bӑ�_"6u��� �j���V	��p�J�`�E x�c����������5?\Ǎ����3L�Ra˟��m���\B�מ��� bW)�����"��$j�9��C�����Ы�������tUʳ���F�
���TJ�?sV���TJ�Q�%�`�U����� �wJ9ͺ��4��
d��L �p,=�V�'�$P�p��"�@��HK�u��܃��0>�O$��bqz��W-j��)����{��t�t�_��YG9�՝�����/r�I98T�/M5z��(7U-T�1�>(6!ДDp���Ǫ˷���Eڵ�3�P�A��c��?݆���iYHH_zS7.�rK����c+F'%o����\{����vM*��m'�6�+3?~�Ḵ��|�.�G�1���-7x As���l�^��]Q����;h�-�Ɖk= ��`�L�o�--�UK���Pr�fWw=����5�gU�=�4��#��f��p��r����Q6jI�����!݊~颢�ۇ�	OH�S�h_���N�r�I@j0R��?ȧ�w��/I�x6ٮ����-��g�ߦ�@��1I6��*���,oo:�ܺyq4)�Ҹ�� �:@��L]�z�X{0�/�r�bL ]��'~�� ��5fS�[B�x��t��`KZ�l�el����I4�S���(Y���[���*BB-��B�B�	U�9h��������7���8�I~d���15Ed��jh$�Vl���Ffȏk�yE��[��3��(7�tx��Δ��	1$gv�ڻ��� a645�wq����-�[�P�l�u\���y)��؛�p�ފ�n�d���0(�v��	*��X/ I�j`8 ���Ը�yÀ�𸱻��UP 	�Uf����o�R">��Йgna!'3SH@@`˞#�ĺ/]<lr}h�ɧ�n��F��8��qzW͢������^E�6Ə������bl����M����Ms�7`Y���/��!hg�S*|[m�nˁ!���D�[ng�DF*��+-i��e���y�p�e�8��k=���5K����P����(6����Ձ[�@��2�$��O` �0්���~���4,XT�m:����@�cc\Fn��
�I�g���MC}��5�飴�:���;48�����ᷫ����{0�{$�B������	�xIl-~��Ƃ��	<���hg5����j�U�M�I��瀯mE�綷�w�����A�U��v��9Z���]^]�377��~|_
<�� ��̟�x;��w2T����SV�Цk��H�:�o���y��-ؑg���ْF�ϓ�����=�Z��jU�E���qza@�C�sP�bh��<�9G!/������|�ɒI��>��R|a�/�ƿeI��$���(y?V�� �ѝ���3���P	��#III���sVByQQ(l?.H�x���4���8B~@�x&���'�Y��<��)g6�bJ���3����]�����l���޽���-""x��v}"π�&
���i� 1R*���#5�x5�?t��b�p��<��MIh�t���n&%���Nh�kpp���k /XY 5䰘r��eβO��xps��l.{�^M��l�* a��� ����؆�`*	�6���]�����»)��I��hwe���0��a�N] ��`*�Enx~v�Rn��tq�kZܧO7q���Y}��9�B�- %����
'��"hց����kPA׬�9 ���{��GG%n箦�u�@�Ά���-���g@��K/gl�Cgl%FaW=�Re�\���q��[��)�|�Ғ7�Mn?Lk6[W]ҫb�iW��; �H$n����7����&=׹#������)���AR�J�RQ�d`UO��r��$�|v�V�o�l4a7܇YoL�i��첮��e�������t� (R������<����h�	���}��%�����N$B��'�ru��L~�q�~�W����^M�g-�H���p�32:
0����X��l;Ɏ��6��V�䝡��\����0�a���y���
*%�����J��I:�
듅 �T��`�ѳ~'Gǝi�GP��g=$�iDq��d>�����I@�w%��Ot��H�8r��<�ċ_e���p�g��̨�u��on�y�L�=mA{]���8�bG|e0o��b�[B�,_�O 1��6��i	uA==��溔):k� �AG_��w��v�e���fgcc�Й0R�Vӣ��#:8��Uez{ߡxЉW�á2�V�w��%ҢU���|ȡ`))z>]�p��G�g}��nb$�{��3�.,X�6:xN��$f�i�xe���]�n,����͖G��P�l��zuQ�:25�R��)�����Eg�����`����������X���ǽ4�^1�1d�z�L��,������+��f�#�0�2S`{jZZ����(�-���3�r<��_��"r�邱n�S�5E9�Őw��K�"I@.J� ��bj+Sp/��:04Tъ��ϰ�72*D���2kW�'�ګ4�zy���V/��ٹ�^ׯ� 409�軄���mO��E=G,.vC�j41K\�2b��+������>���T���P}���%Q,Y
b�R��Ԕ�����cPSȶdX��c�o�Ru3�b?άB��'UIߥ��p�w�˶F�}!�2^>\�Eh����Y9�<	 _������ͣc��BN/>��سW17�����srrv��pȘ�+���)&<z���c��6n����
�����QXA`@A`W	i�	EB�;T�:TXBPR�s�!D��a:��� ~�g�����}�=�\+��k�G@�Y���u��Nn9�]s�yGA�2�vonA���|��rF(���}�!��'l�rm�B&��+f�2 E�{q��&��ۋ~Mj�o˺?WX�@7��q3��V�� ����������Vj���@��
b�c��+<@-�m�Ėp�N4H�y*T�.d|6���
V:���nn+_H�\��q���\*;�E�C��w���?5c*���� ��ǧM+|@@ �/y-���M�Ha��"�;��	;�v��o� bf3�!�/�v
�liyB+�k�cU � %�4��q�S������5$$$;�#���k����?䈖|	��q��y���Þ T�7�	���r[��$lb�S6��5�.y�t��1���D �M����9tV��osW�w�.w.{=�(٢�_��@k�[�B���q*��x|tJMC���Bm���ZF�V��#�k	2�3����XĹ/He�t�(9C~Z��i>����� ���x����� �iB�e��$�����\�q���+��sN���{?�%+��)�_b�ٸkW���j:/�+(��!K�ń>�=��%6��0���a��&��~��Ϝڿ�� � ��۫����'��?� 1Z�*���I
?�؏��(ԭ�.�p	~~��z8���S�:�Uq]���^���G��+�S��ώ��&�WhY��=~��rs)�����u��hu�+�s-`'�.h"�%��W�T
��E�F�N��OGЉB��I��$e��П�$��dU��ma�%���@��͸�{M2��CPm�[M��){g�h�i��W��Q��@�:.qtT��TL���=vJ�_)�k.w/#d�s��Ma?	b�Y�dr`|�-��%q@�@9��kf�h����o�=�g:\�Z����Q����]ETW=ڔ����㺘%%��珃]o���|�<+/�����eQz��㛞~�ƃH�˵��<�Q	�ѷ�Ԟ9�-�U�='&��9� |�@՟ W����p�E�=�vhv�Tj,�ݏ�'dA���A_�S�c��Rt���g�UH�I��e�fݔ�h4�ȿ��@"
�B�+1��_�I],Fh�bq����
������zßI�HC�!��.ۋ�c��\��YH�ɵ�R� �#n������[���&C;�����mAپ#1��ֲ�k@fj+ЍѤ\�c3�V  Y�5��;���;� %�\~e�U�[�x��Y	(�����}y{�ѫ���n�[��9� R�l��FF�ம�a%F�z��3���sF�<׫,���
�(����+-��/Ҏ�|�/Kc_ov;��ڛpӧ��|`��h3E#^�ͤ��\��_��m��azt���.]2���t缴�mj��x^��QHL��(}q�UD��x�ɳe��(�yG�޾��N���_!���$0 nO~��ް.U���� m��/]��q���Ȭ����Xf�X�,�Zl�[		�\����>��S��Ijkkc����N%��������K{�(i�2_��x��ˮ���Ίt��u���|Hq,M�.Ӛ�9������� *xK䤜S�)Ub7V���a3�D�A��X����˨ͫ׷��ѝQ�ݓ���J@6�AOx&˿�#Mf�9!��yu��-��E󮯭�9��(����~	6\�k�'ٗ"� ���fs��V�8�t����l������<ɻ�CVj%SXQQQ3����|'�ml5<t�_��N|��YZO���������-��kЊtY��jeffR���\�J�h�W��̭K_`�\m���Ye�� �0 X���h��B�~�����\�r*�W�QW�܎'I����}��m���'�vdm�f(����J� lY ���j4�k���Bh��\�|>F�K���v�*��W�Dڗ`��5W�{�����ņ�"�����;{{qU�_����W��h��+3E���%tW�Tb1���k��#������_.���A~�����z}��io�y]N�OV2z+V�%�M�,�9�sM���A 
�� 	�~�֠8�6---N��Vkv�X�p	�s�K��U�$��⻯�6�.e N�����"%%-��.����T������\vz�!� h�Qh{��k�ϵ�˲y���� ��jۜ����u�������*�""����Ȏo^,8!��1r����5W��U�6 [Z��������Kz6QB6n+ ��#��ҫ6w(_��G���t5�7X-_��PWW7K�N;Z�&��>�>�\ᙙC�M��p��D�����-��i:�}�����k׮up_+2D�,?����c��D�hlUdd���Oz���*�@��U-�A}�SL�/$�멧�G�&���J9��ը�����mY��|e��쬠�b�< _�F����o�g����7���'�m���҅�O27�j�xԩ��>�U�X 6g��U���t=�-' P��ҫ:��.�~���U�΢,��������..���{��/���N�^�_@ @������<|iܘ�s����0�TĀ3̎��/�|�{-��w�Հ���XŚ��ug��nL0�j�/:���h|7"���ٝ�:θ������T؛.a7|��*�^jD��of"{�h��O����VV� �궯A��?������3Dw��(�R񸸸䥧��8��kP�?�7C=9����~
��: �u���|�-��}�A�e�!�<��0�� ����:Sⵉے�r�ܧ.����rv����{�����sN���[�l�G�tc��c����'��
Pe�jM<�ʣ��R�i��6]�}h�"m��T1
m�d�;�������L����}���tͫ)��.=�~2���) �k���Jn=�/(�K	-���o�Tf5��,�S&��a|~˻�B�7%C�4Í�P.5p��&$�g��UX}||��
�Dv.���C��===�8e�J)�P������f��Ѥ�b�ԍ
�q��_D��əW��m�����ӥ`������,3�'�Xb��9K\�I�����M=�A^����}�<�c��� �C�\zE�����Xj����=|����?K��
C�B�/��3Z����x�V� �%�����h�P5���ik�4+�2@@-��X��;!l�#���#?~���h�?`YF�����L��xN/Z.j�[�W��rF�ŭ�|nx�^R:m�,�U:s��̘�Xx=�����Gx�w�������u���bK=���/�m�T��8NC57����1>ᮁ��eu��\���>���>�ap�tw܁�,Tx|�\�¾}u��P��u444������`D[��;��t��C�;k��Ĭ�i.ĥ��-���@��l����g��Қv�#a�%~P��}%��>�NQ���o�'�O�p}mL�̶ۘ*r������u���PϬ��$��mƞ��� co__AnnЯp~(��{�6ŏ�Z܁�(e�$c��g���;p����b�0��@ 	խ�g]N%����i-[K��ד{ע��Mx��mu1��]���"+�"��O��:�<V��"�R%��yg�EJyUs���yd�t�ߜ��x�ĺ	q���kM�L4��[�STȳ{Z2����Rq�&+Az��������e�~.{��� �t?��ث������]o�
��,�Ғ�D�/@�b�W�ӟ��l��~E�C5[��c,�������F����ކ��������{�m��
x��M��e�k][�Y
L��rG�����w�~�1�X���8���<�~�XSǍQ4-�BlO���N�!H<�f7n2��X>1!�+����C��	�6���������* �%�iR� ���xyy��=(?j|���.�N9��g)��bn��?�A�dr�M|��n$�8� ¡��Zx�[Zק���]����C=�Xm@�L�
�g��t!�J��e�_���y���3I�� #,�
@@-3�����Q�ە9���bb���,�5�i���M28/���Tm�=通����&��<��pjq1��H�J��UXZʝ�����p���~s@3E:w���n\��C�߽3�Ϡ�D�vܾ�C�x���A!�ӆ��Dy��Z���l������l�ΝV��;`9Y{V�D��
�	�FZ��yb�h�{��4�(���M�~�����)@ 䓓��ի�� ��6M����	���O����j�?~|

���
 rc3��S r�B���1%h��{{�r��>���z����F2�w튑��@��$�|�q�������4&�SC�V��l�p<��ؾ��Rf|�Z���9�eu�b���d�~y���P��`�A3ʹч� �M+b ������D��y��U�ۏ���koEў��Be�y1�����=�Z���@���(�GXT�ֻ<_�K���$����S�
��b}����P������)���N�f{�s��
����6�-�V�	�{�`R�X�3���Կ*��s��i�'�r�T�a���W�u��j����s��RTVnn�H׸���s�j?����tܦˤ�'��9Щ3�.iz�ȓ���R��K��W�=���t�;r�A�΀�؜��5yd��w���9e�'�$��,�������r���ӭX'�T6����W�K�~�մ⹁)��m�MFG���"�{	�c��!��/�	����|�_�,lY�u�Pf�+j+E��ת�G؍il2YGCmB&6I��뉩1 ��f�bs�G2�	��Ƭ�E����TU<���^ ��kL[��w�CO�<	hȮ�r����p��@%��5$����Pg&�R�R��Ï�L5pGM�>X\Q�l��cW�k~���9�-Z.{xd�"�|��
L�`� JB�E755�ހ�nUp�s��D�L��I��zL�h�q�~ )���E�?@��	�
�ק�0���/0����Ⱦ��a���\S��Ʉщ��Z_�|�R��^�g+���a���o����mf���q\�Ts����������t|Fcͪ�55��FC���G�Xo��(yJ �1���IɃɳ��~'a���������	��p�M�r�` ��E�T%������,�gE'ם����
�@�p}ڴ����g��-��d:|m�'{	F⟧�jj��vZ���45}D���2y*��G*N��HFF�Y�%�d0҂���ϗ��m�lVE6�I��<���A���#����~LC��ag ?�mG3@̳����7cK����&�J�G!Ղ6�RdVJ�͟��-�7F�,��J���r��ϊ���������\���4��K���Ю>>���;+�V=)��B�bC$�0
�������)`�Y[���T�*b~;�;�ד*����o�#��A jU��˿�h��E`c�y��݃����\���rp(Yu��3�{�4�@� ���o�P߹S7��~?:��v98��"�������;	h��?�ʎ�؛= ɺ���i?���:�S�V�_�����b���\MP�X�ho���	��ӜS�� ����wG0r�sPx��~J�����+i�Ny�C������A�{��6���m�@WAe��So�n]#d�P�Kp�t6zx��>��R���J�y��H,�{Ǟ�d&�9�Q��hM|[�p�ЧBwsZha*�mmm����r���R#.v�sѧ��T�0�� ��ŮM�e��Z���]�J�~NuI��������&'��O�]#�b���eu�GZ���K/� ���f.��چ1�V�t��%�����#�q���>.����#i�V� R�K�~zP�t�Bsj���Qs�ՙ�D����gb�zz+-	q t8��<c������%당����_�jr7�O��
�ܘ��m6�t���0�"�� �g4�!DeƉo���u�������%��m�;�iil�>^`ޚ_��C�0IZ�u!��ֶ��6�뾚�.��U�k�BJq�	�,	�����>jض�F� �Mջ,�SMZ��K"ƃ?��U�"Ϊ���f=�Feo�]� o�T,ܱ����8�|�|�s�s �l�nE�;���=��-㍫P�����4}���V����!�N�ZG�CϪ�)��q�A=tWo����0)5F�j��^�k�/�N��A��6|y?�}��.���]3g+��I!��G� ���d߄��& 2�d�/���}���3<5�Nq�=Q%Xw7�8�ٛ�w�և���O��6�
��04���oBB��	hiE:��_Q��ʑ�W�Dj&=�W�%���q�2���ߡD�9G!9�2B7�D1#EW(���~�� #2T�o�	܅�
���M9��!򖆏���I@^�S�ݏJ�Ee��M2��7DT��A3���հ���P�/q �`�����to�\7���:r�aKDUom-�tM��rk�̖��:L%����
 ���'��'rF��/���u��Gwɤ�]7l���zyii��A:& �ol|\^ ���}[������/��PNz�'�<@	�p��/���]�:C	p �c��GCn6����~�v���xI//��|e9`��A�P�j�q�Q�R� �����%6�s��gz���\>�txP>'��	D�4yy���cW`*���ꛞ�w.�oI��TP�=���h��Z�D�tYHA �J���*_��Y����#j��'M�->c����m���V�����G��H��Zh5ED
z��м��˽����e�e��ֻ�%�$�2����2W��&3J�CɇP�E2Z�,��TBR��uIWO��S<�������ff���wP+���ܷ��&�����s�,�����2y��w-�x���W� �]�q߆���jƋ�5y#;����o��X�_&$$,����0��o��jV�ag��@��5�[�
��><q�D6"5�$S[ .�ᭂz&�T��o'l3~���$���R.�����XĽ	�T(S�?�j���'��!"��>����~���:9�'��о�u~�*��[������]k0➜��{B���
9J�"ǫ�����Z�����.�w��+j?0�ΰ��o�@P��|VΠ)��p�ky���r��wtxSխWW��]���X���r�mm	@�QA)��Gc�J�#W{���~ǸC��&��'n�8�����U�8����-�"r-�{��׾��&��៖�gҬ���r�nvY�����';h�=�GYZ��Ą5�D��$ "	Ll�J�����E�
b\^�:�n:������Q��笢���=��N�i��33��z�>�ی,����,)w���2Be���;�_���@�^s]���dӿ��W�t	or�%��C=�(���q[��蟩p�o�C�lBb���Xf�%(*(@�����m)	h2� Iy������l+�"�گj.O���ꏡ��S��/<�S^ {�l�U�p��i9�^;a�#����I�����*���F	 -��1���;y�c�Q- zɧU2|�5�1����� X�&%%]��G�-{������m4]!����R2<�_���dQ/-�$	����+ ����:89�ػ��� ���ɛUu��h���2ޛ)x�7��4v�C��������!�?ۡ��3��v+���\wu@��N7"V�|��Q(�u\OR�t�IB��Yf��0�"��?��$P `�Ag�7Jo����I(���B��V/�	%����>R����E�6Q?#n��T)�o����|��1Ҷ(��6���*�sobW	�c�*�^�ܣ�3���e�<'p���aM?����bW^l���#���3�S�7�{M�ԏ��݉~{U�Pϕ�V��n�0G�ޞ��C০�{����:���5�`�K�Fj�>�])�n5��p8��/������%6�* -w֣���,DS�x�+.�G��E�w M�W��e�MJ��Q���.�(�E��w��ם��!�����-�����	hy���l�;n'�_`nN��ןN�6(���GD�<�K("j�_ ����W�;�ƅ���7�|u��u�5W*d�VπTw-1&S�p5�P���ӣ�Z%0�>e֓�?���ho]�+ ���/��AOJJJd� v�8�D�JN+��[Xu����9[U7'�g�.��&܀'�h(��_��|r�б8m'p�T��=s��,=/�M�<>@m,i9e-�l�F��ĥj�`���Z�;�]���dVc�L	��W���H���C�\��˳�#'��s��y=�+zQ�zg��\�/	�f�s!�}8�o���Z�Ǧ��<]�u7S�s_��'���O.���եde̬sv��eX?��/OZ[閨�ϴUWd��8SD����(�Y9W�ڡ�h�����
�8�\s��Qy�����dd^^�pZX�hyOr2m�.n��}�Qv{�Y�X�ʆ	��o���h�r��:����_%hԕ*On:�X��I��^���+B���8�Z߂��ƴ�J΂�u&aq��s�!��z�(���^���4����\:P�R���W>��y�/��6j�ebbR>�f��Ps~�Tj9�~5��(:�N�����ӡ菟b?~�Z޼��D�Ip��bi�N�"$��߼�l�s[h����>������TP���[�b�4]���X̄�ƠG��vla_զ��y߇�'4.E���?���m��.��ژ����*�z�N�(�����c&Q�l��9�:Z��&KT~T��1�u�f��|c���P
�-�������+�=vJ��c,���dTT���	<�cy�W�R^���yj�0^b&¥3դ���\��p�YpEPh�q�6�NQz���*���&�#>11{xV�CQQ�������On��#,L��������"���´���|[r)���������=Wk��s�|�䭭�X��Ӡ��96ぶ�4���~���s����)���1t����Q�t袰�>>��呷�/�/{>�B���s\8��gs؏gR�3m7,�)�F�\��?���i=�5X� �3� ���Ne:
�/�m�Th�4���fN�	����E �/h�nz�{^�7��߿_?�!<����ޥ<j�}����NY�'C��������<Z7��>A��yz+D]����9
������";B�~M�Q>�G-�5��R"��W��7AǦ!����<��}�,��g|��'|�V3���o�i��n_o$~��5��"����ji�ٸI7g���_� W3�`~ۙ��?��B/���Y ��a|�XW�݊T�3��<C@�R�s+mGyD�V+���s��;'#�����{��/����˨F�\RRצv��h�Ǿf�--,�`n�`fR3>�2����A�+47*���՗��Y�L���j�N�,���{A\/������b��}��Z
�&�u�� �ֵ�����1G*)+#���L��X����}<�Urn�͈p�pu,�sy�VXdW�L�p���&�����t/Ĉ<��!�W�41��h�z�tX����	i'i&R��Y����h�>O$n��)ؕ��[3�jg!*��د�/�@�w�G���7�.8���	'U��ї�46��7K~�[��.����ؐeP�f���	����(U׬;����潴����}����4�'<%ic����/R|��K�[�/��2�4�%������t�?�-���֠v��2��ٵ��Ղ�C�yg����Y6l�#خP>��yT���V4�k�y�4g&$5G1��ѷ����d�E��a:� ��?�Xo.�8���9�M�z�D���e��NP�Q���W(�0'>.��į�SJ揮/=91�/tO�E���#GU�J'� zk�A�}�߸|?jz�����z�1GFFf`ż�{��i\��R��Pl:=@D�����k���/�~5u�N����V�T�;���4�=�/?�3>�.Xj4~�ߌ�"�L����	#v�a,zsb}���9���Q�e�JE-���1����u�|_��3�֠����������	�6�$�?I���]��+���|��u{8�����K�T_�(�fM��ҋ2'�d-l*����Χ��WJ���ti���1�<����(jV[G7��m�t����o�(�<��9ڵ�nh�ʏNAn=��ޕA^�Dlu��"�i��F��j�~�3��|ւhKu���(Y	:os�3�5���\؂�$mr~��I��u~N)�ҳ�I=�Z�O�7�R��I)��/���b	�+�M�����xѫ�X�,?����ou���LB��Y ��ݳ<f�8y����L�*�	a�fqY��fh��kUII�'Cǃos���?X��{�"r���\�e��	�sݴ�ŏ[�d2,R<�O�MҒ�������t2F%{'�����Y5Y^\|p��7u�3�鿯rw�� �)�����.�?���,�����DD_�����CR��E��b�w��ق�eZ����Q�Yff&tpxtT�q#�Y�
�M�����s���<�{]�)H�hyK�[=���6�]����y�lyg>��:�|-.<C�%,����t����^��E�I�R���49�,�xd�bO_Bo�e�@Y�@�;J���}^��@�J�i1��^_,F�i���Z�i_c`�Q�`��i�(��參@\k���QZ֩���Li��]�{dx���<ϔ?�%�ޘ�������9�Gd��	b�e�A�s�{���(�NN��{y�(�a~nnGu�g�J�P�����[�)�߆��U����3/MӒ����C�yQ���)0���I�b\˶�*:����KxXB�a%�BJ��NS��V��} �R��j78�(4��`Ek�0���Q��l���{E,�Xv�v�9����[	����u����:~����-�e��V� �5�9G!��:�R�o��l�_OT�:��+����Է?a0�
��b�`���
a�������:�b`Cd�A�L'LQ�E��	9���+Dr��=��[&Vv(i�2�a��rL��6�I�v�}*����V�s���h�S�W��q.�	9
�!�iH�u�wƵ@S6���G"C��#H'�G�U�9\�Z*D�`�:ۯ�z �M��ٝ{�K��RXZ��UzkQt���X�����,�|���K�[��N���cKt���Y��
L��R��A�uO{�k�ʁ����d:O
�9^g��6����0~�}�I��$�����Q��5OvBGQ(I��""'7W�\vF.����xſ��ۡ���&�`��~���~K����?��3�IN^,u�Dz,0��2(�ĩ.if�=��e��F�?.���J:���o��BTkP��}#�lOLa�w�����p�<�	��31''���gW�>��9�4l�6W�PX��_�et�)T]�?.%'P~z�cdd$ݾw��y�s�+��n��6�����Q�9hP3���� �����J��D{ �s�;�A�K���Ax�Ό����{Ή����Z4NCV_귨�%����	���xG[FC�-�����6������"� ��	&�������������U��!��qv~��b�#z�l�����p�n�,;�߹ j40���c�70X}�E��T��vy��+q�t|0��L |�W�/t�� �ݴ�D�20���t��þþ��F������0�#�r��;��F�&��'�����^�]�a��U�H cGb�_�R��]5u��w����#�宓��f�C�|���/��s;�;#���L/?��G������`�/	��8�x�V��%� ���mv~x=�C�$��4bh�b$~�ޜ&Ee��`*���9�B�:�9�^{ˋ��e��V	��&�\(��k�"u'���u~F����꿚/��Ө4w��]�rV����JB��j]F!�����;VW�T݁Հ��!#d���?�����ӢGK�x��l�x�FX�<��i�3�#�yx2pZ�y���P�*p>�w�N5�z>�%CM��GGu���Z���
ݍ}y*��i&*Fw2(�[ֵ95翉{4��\w�w�牊3��z*��ӄ��۔!�$���fuN����ca����lJ����C��+������C�"č*}�Ӏ����������uq��)m�a��/�jg���j]� _����dq;��B�D����J�ˑ�]K�]� ��Bi�D�.�;�����vK��7���>=§��Qc�^�i( 3���5>��1!��m���׏��KU^)B�y�
A�\���.�Q�+���F˳������,Ӏ�`��ո�/_�Q
�J�~�\����Q��]|<`ݯ�a6���3��G��~�$ϔ'_���u	:)�^�Y��x��We<뮾��jE{��>�.���K���5R�Ni�����d/uz�7�=M�'0j6��oE��փ�f�r�؟?K!��`�~�m	OB�N6��/����=���Lu	&�Sz��w	�M�Y+sQ���Q7�b���)��x�$%��<���V\r��po`غ\]���bk�ͱ�Զv6�{�X�ɹF��k��4��t!#�tlw{�enș'/M��JH&@��%o�|�9�1�
�Ha�m򡦦.X�[��8Cgĸ��;�G����4ΘMIB�+��jօ�������te�"�� �ʔj����s e��5C���~�����9h5�x�M�F���>!7T�^��/&�N�e��$�|�q+,��?p8<�__��p�/4Iȁ�82e" �c_����@Y��t@p�$ә2�, ���N�J��YXU�|�4|���B��BÑ�����PV��tr�����,�
�9Q�lY�õ	�6��)���B'f�$�_Pa�4����f��ù�oX�h��[��v��]B�JP� ��"�*CθX}�ꃗ��o��w���٨�^g��B"�6T�;��t>5_���r	 wyΘǿ��%&"0�@�c
k���쫸\~	�<�0���a�'���3����_i�N���o��g�X4(��+�!�YM8���`ζZ?��'YEst���ѕ���9���+�ش��P!���6���EF���H���~M��*�p8tt|��@��^�wh"���tJop�*YN)���4oF��ΰM-���O3�`kF}9B-L:���'BX�5�S2i���}�\L�ŵ���6�2Gկ��}�J��^p�P�A��Q��`�{���*W�v	|��F$v���Ȧ��^���f_��VBk�T-��h�Vq[�0������ ����[z#c@�G�ǽ���d<Vˏ���۷���]G�0�D��*ӎ�/O����:�=sa����%u��(����~:���p�x�
���**�!�
�m��d[��[����'@x�>vW!"���
_�GF;�њ�6��>;w��kw6BP����M^��bXM�p���f��I{8K�KƹW�	9��GvP"`W5��p�p��y�M���+\@=�>a�6����.}�eX���%ӭ���Ac-����/�qo}[�̸�&\zV�Re���f%�k@����^p����E�7��2�M�}�)/B������w��{�>�ӓTh�=�mR��nge&������o������!@��pu'�|�-�w�r"�,6�
���^��{��	{ƨ�/�?[W�*W�*��(�P�:d��?!�� U�p�?��3?*A#$������������5���㓅Z�����]�=l4~�ݔ�/���⮮���ץ��SL��Д����	��<\���%���4Ȩ��`�/v�U��\����~�0���������S���4���W g���eW���G�W���+7ズn.������<�į��-*��rg<_:�:;�L@�����9�`������U:�u�L~�u*N���������x�Q�ή��#^��u}}QΜ�+|��z M�u]w)����9^�� �hɂF
u�G�|||��YlH��P��&֚qßU�UW$���u�=�3�1��h�R����@\{��gʾv��.���D��V���B��W�Q�S]@򟟐�J�G�<��&���6��Fю6 sU� ͣ<�3a�a+ U�E�̴^%%'G��w�h�Y�R�&&&���P� ˂�&���L�uN%�ӳa	��=�=l"^[2�ΣD,ഏ�Kh0��z*.#������DН���8D�Vsue�b���meC<zn��������B }?74�7Л�J}L���1B��H��8tw��o`�V@�����WBэ֛P���v�\�84���#ګ,��*���8R�O�9�{�;P��{��Sl��q���v×�5e#_�(/,"ҭ�fn.��>~� "=�(���X�:5�����4 �)Ӵ�����H��w��nŋ���dʙ��}�E��Jko��Zr	��$ ��Bm�����e��NC.���v��I���ț������W2|��n�,��������%�UPm�< ��K���r�j���[�Yʏ ] �vwיv��,���I���I�i�O�|�j<��^1�Ku�A��.s7�̌�q��$&nT��8R��b9 �	�:;%�vQ��i�o�T#�9
Z!Ǵ�ܲ>��%έ�o<;�����f�8iy�W���ᖂ���T�T�f��+Q�U*�����t�:@�#���W!�Ζ���X;��-����:��hHd���k�3��S��N�ﴂ��*�ȿl
�Z�r�G;����q3��������������o��v>Eu�x7ǚe��}m)��E3�9Ң��ͯ�Q������ps��?6�>PfVJ�������X3nO*а�r�CM�5�zB$,tsk&��'��8����G8���*uh�_ٺ�&����}�6m|�Y߃*tQ�{�Nrv�"�3�!%#���)�I����6�.�,Q�&^�-������̙��Xe���lk��==k	))#����K���m�SD�q���՞omgg�k�No�:�@�˂%e}��->|	��i_Ӎ�С��6��H��о�|$�8M\MA[����x��G��@��E}T�-�Nq �w�3F���<K������)1^��A5='~dA���2o��&��ع$is��<|F$911a��k�B��c�T����!�JHDD��0����d�z�/>��%���$F�k؀�� �+?x�m��ۂ�x}��{�tW���j�C�Ru��/��?�!������x�B@� �����mZF��j�&���S5j�X"����Hڻ�^6Ϻ�������$g����at�i��}�UTF�(� �@��`��]�q;U����B��{�����i����ǖ���{�Q_̣x�߬��>e�*'���΁�ׯ�?���fK�ק�
���GE[f����$������J@'#t��OKLhDj�Ԙ��XxS�ax'R����Bw ��w5hF��=&��ݬ !	��5er�	�H���>�H�2��\�\��	,Oη�9ǁ�+��~�8�DT�T����]N��p�+d-z���P��)�;�GNNN>�4�];�c7��O�������6B�B�|���Ϝ?�bl��L���g֏��R���^9M��Q��I�uKV�o�+	�2����u�����E�U�udј\yg=�Z�k�l���pS����[�l��,��i���_�������Ϙ	Q��
�����<��|�4�S�׏.q/.-��a�I��5�R^�09�	

rX����mf��=����-6.~��:[�GM��n�.dV:���談6^(_�A�7w؛��7��%��V~�P�э|��a\2��M�M�v-�WՖS;{�GM�-	U��0�Ǐ�S��n޼	��kr��>���ܕ�o�����|��nC����q^-�x��?�F B�-��ݰ�.�,dH�+J!-#C�r0鵞o�)R.ho��1��(Ǚ�D��	q���s7/�=X�pf���Y�CE��g_�n������j"w	f�-��|r���,�}wL��O�6.Tn"�|�J��ի��_��Lk/
nŽ�����ucœ���xz� ��tu ��|{5��],���[�SL�Q�,��R��*�z�m���w�E����m
9������O�H@5���� ��&
�K��eX9_� �-
$t�I����]Y��5�MP�
�E=��{�n�8��Y�C�^���ww�e4��bz�'��%�+�`ħv<)���eW����=�g��ym�>)��$����faa�{����Z{���p����.���/vTX�* �m�����ָ�\�M��>'�eJz::y��@�Px���/.��$�>���t1%��k�9X�J�H�Z?�+��^9�{� Z.F�J1^юS�V�������?br��3���b����ZՇX]�GF�BG�᫈Ɗ�e�v=����9S^U��G	�D����1������f$.�L�G��,]LO__n�]&����\,\p0[KYc�����;�k�a�U��egg2[)����w4BK[Z��x�:�\�ة�_9�V&�Wz�� �?e#�ۼ�W�}���dffV�Y�A���1�$�eg ����s������;䷉�)�2>�O������L	)�We��ލ_�~o}z9K*5�2����>%f{���Û�C��C�:�89t�99i�x�j|Β+��
 &��^��s|T�7�sX��ܷtt�䫕,W�,����) l�t�X&S��:f�������>����{3v�5�:* �l; �y�) S�����$ԃ���2�����u����T�j\Y�r>�n8���N`��Gj�K��v����~#?~|R˿u⬣ma�p���8��!�4F' �n��}�T�1.�L+��o�aWLED����Ǯځ�		I�zh������+b��{/b'ȚڟK+�:\�Pܐ߃�B�c\��K�Q0�~�(��a�5f[�IG��2"��knm4�l�K�5&�b_kO���j�ʁGӊzj\@\b�������8B-�����~0����sg�pZ��_߰���IM�
�m��v���"\d��!��2�*Bv����lb'��4���0�[�z�/m���]�q��|S ����MB<�m���+<�w�������ٶ�`��n u��l��ӿ ��!7��q#`�ç-��w��;�g�G'��B�V>ՠ
ɯ]����rB�33�Q�!�]��7���-�{{	).�^ϙ��{�o�q <� �İiC��|��<h�~q��)��]��lx�?���Y��2sD��A�e�Zy4Q��@D�R:���d�z-r��|��̎ҟ:U�(�}��<�>vs3M�p�#/��sKˎ]=�b�2�a�����V������gcu��zU�fvĝ�!��� ��k��Ŝ	���_2�X��[oF�4��e���W�{�5��ƨ�?2���7��dY��K�\�U�?	��WW+�=ob�4�M�� ���N�i�e�g�#��z�U�D�%�2dXO��l4�pl7qSP��j����֭�o�p�R���zR6f_l �ӫ����� ���pO��]�T��8��#�"��j�q�'G�f��+8�u�ʘ�ړF��0aaaK^�J�d��TSid�p���޾���SzZ�M�$�j8����Hz�b�+Ā�x����k�����hxbb��.j5��Ғ�SU�UĿ��`X5��oߤjL �U�}����N�$d��u�aMfM;ꂫ���"��T�w\Q@zG�J/�C��"������^B���C@D�I	�tBB����~�%?�}w�9���}�s��H�UKo&�e�Ϟl�}���l& $T����e�TY��������9�Qd�̯�GTp����(C�\:���Qz�q��\�cy���ّ;����ؼ�����%��	:,|��'��CoK�)��pD�j|�#J���jq�:���[gQ�_\RRQ\www�&����2~E��^]`��!i�����2Gޓ�f���$�g啕�_�̅�ea�����a���_ �XI��]�u.�^V��[�o�QÄn"�I�}��N�1�� 7�Ã��l����nTʲ1�%�j���Y$0z��_#\�cC#��H���eM(M�0����zJX5�w��s�'L��ҏ����4�D0���p�Q��@l'	H���R�ԢJ��o��q�0*+ݒ2�!i�$ͼ���t���/D �Rew�.�+�>(�����'��t?;���\�����E��z��bf�߹�08j3v����� �CxWb\gIH%�{y��N�XD�o_�~�<}�9�{������kc�9p ��N�$�J�sC �4;;`��,��q&{����z�<]䔑����;�����t�E�Y���P�SE��ڽ�ܞƋ���,��O��ݝj%�j��:C 5��p���7�VҠ�L�a�&&S����j�T'n͜{�\�����hZHXg~f��hg{{�����I�f۠^��h�-��`I�LC�s�� n-d߄��T���]pdI�|\��N�&/`���_~<���~o[��ۊ
>|�sV�E�w�τ�uL�?}M�Do��:���D�9�������ꇠ���I�����|
�K`2{��N!�@����;�T:��..�����Md��y"�G>跷�2�ʋ�+볲��%j����c(�1W9���>���������p�����vN��Q�h�����67���0���Oa|#Y߆XܥV�3�4wE?��;�QMoo��^G�pIn�_�*X��;T� ��A7����
� �C��"���3g/.�d�Ũ�� �87��ep�b�&���r�^����/kNtWF������rkRcufZ��c}���[�+�g;⅄�r �Vxs�Hw��P�\7q�o#�jܳ3�V4�F��6sA)��bêvA�*�b#�&V�����e�D�4�"}Sά�_4:F۴s�j�d[ĝ/������>4My}wf���9��4��Ѩ�����c߾D}����xM����Pa��-at@�gyJ�\8G߂��1�o:�v������u��|��/Guս�S�$�aĒ���b��B�ޞ�~�p��p�J���;]]]�׽K�|fq�~�b�Ĭ�D�N=y�~R@��{
�H)%%��� �wG ky�HɌ�õg+9�"?߮�ʂ�˘:DY��#�a*O�Id|v�Ī�q>r�U^�Y}zNEU� /O��<Z����k��p�L*_܇�![�����i�I 	�a�gΎ��4�0 A֛�Q�WI�-qƾ�&��w!�8����5~D�4�*[�NS�)r����z�Ɗm��g�aLӑ4\��;���N+s�� f&&'������G�^jz�.+����mY.dGgu���!��Ë��o@�r���Yn�^�}��_�v��U��$K:C<��nZ7�ҴP�g����\�Ipț����-$h������� ZS�W��oit6�9��4���;X�N��ϷsrR�R�])���\M��a,��c�eQ��9pt��p�k&%w��yڽ��謫���ۜ	5eX�߄cll�r���AqBJ� ԥ$��*D#��?�u	@�(c�I�J��e�����S��q�5�{B	-EA���'��G�l�O�=mH��U��G�K>���a��@`u~�n����\-�k{�o[�4;��fu=?k����l'|7T���Π�����Tϟ�f7���2n��˵0kkP�'��2���&�`��uP|�Sv�a�`��]�3u,�ք�@��\�� ��2t�w-l�lncn���d��4?p�Ls�C��s�!YK�ok�WC~���Csq���g������`f�郌4ws��EX'»L��ߒV�n�C�)XE(�)����e��nU<����n���ɯ�$�-���UiUQ&h@�o<�B�eEmzU��JRB���`	7�N�_;Xa��8˲�#�1X�]��LP��z�/���e�r�I:��Xݗ�qPe(+y5j��-q��]���Ď�Y�d�G���
��56M��}�g�pU��B1t��&M���O��t��e��/0X��\�:�!�"&,-(�8g�j�V '?�u;�����+�1�݁������i(��w��V���u�G�,�+�#������Α��ϑtk���j�)))��46F�cu�ɇ^��݅��1_=�������5_)��p�]���7`���V.���dv�޷�P�(]�}J���IIZ����i6a��. �����*�������a �����������%��ס|,��ϖ�ĄI��������e�>��	�i����ЪR���4|�h��
�ņ�}/�z��@�P���4����!�Xd1`Кyʩ���pY,!h$�����A�w��Vby'�U����g�{L.y�����H"4�%�����ydVV�����-�<��:C(bG,�ߣt��4$R�jj��C�(��Ih*�Χ�����\��bKb;��B\o����q����8�$�p�Mi�Aԋ�Bac=Ϋ9}6�m�7���["��2c�.\\\#�pC"E�6�=)���~����+p��kY�����<��@V���["�uj���R�V̉�x���+.4�vd�-���5��L=n^"B����GFB�� ڌ��54�T����<"�`����⧅z����?��W�SN�<i����Q�xr�D���>E�Gj:��Q��l��ɭ~-�rhI��L����N;�A�ѳ��8}������h�{u�gaN���A`ͳ�J��ޗ�TƵh��i��X�(�#�s�E�-CwP_u\�1�YTz�Mq<����/��n���>A��p̈́�;�++g;�(w��Gி��ϧ}����Bj�Wb�3w�}Ԡ�Y6!����mK��
���1�(:�3��J�b���t��b���3��XIUG�������~lnV���`�wQ�B�if]�h�~/���D�i̴��f��>�Ӌ�`˄
�|Sw2V�����x�Ӗ�F	]}iV�ۿ�X]xS�g/�<˚��nM�
3Bl�`�w	����
5Y}�h�sX��8@��P=��׍�v@ެ	�8,i߾�H�=^s;%����k
�}�Tu!\jw��%���0��u�]g�d���	`9W�w5�NzgQE���Ź�$C���N7��rz�BmH��q'zdS[��i�
����q''i�G9�����<��ı�\.eN�r��X�W�V�.i|Em�#���c�ӵ9��^��)�)��[��V�� �rP*�Ø� _����"��^���lo8(���K�����6�f������/�2|���D~��>�Xw�/�8üߟe�p���=�*�%(-�����궐 �V�,��bF��`�GDK�ߧ�jN�����>��l���åB���1�u���6�6!/ �_�gB	�\�3����źBbbP.?`ٌ Tmh�d�"z�F�3����ln�i����o2��'l����߯=&�ӧ������2(��.
}%L�<��u�a7�n���y��ꆧ$b#X�
�ߚ����<���([�<�+�s�������s��_�h�Tt�D�K����*���*���@�	�6���R���k��O�D����C���J��l��:<\�\e3ۑe�AX��Zf
��93sss�q0N����"�	Y�U����7��i�W)�������0Tj�D  py~�#����G<�ħ��e7�m��{k-�|2l�,�`�Y۴�zTqLk�p�G(�$���4n��3(w�E�5�}��ٚ���q	����MC�0F��Z�ow��A�۴@3��QZ��	d�=�FE]z���v�=w�� �رmB�Y9y���P=_&�j�P�������*s��W%S��R���uwG[�}5J���� �ѣ4� ��v8��� ɺ����\d����Uw����GeJ� �(h����TNS��R��%��Z����A14<�J�ރ�K�>��vZ7�S�}im�g���o�ӣoxE�z(/Dz��#���ɸ�������Z�J���?v"j��(��,�*�<�τ�R�7I�v�1�>:BͩJy�m�.�vԿp��[%���AC�Ž�4=@��_w���X��W�$��ckҀg��c����ts�?�RT�q�lT~?��p*=���w	�x��R�s������e�U'�@�]ϴ��$�"��[#���w^��<�ӀQ*��bXz}��ߍR�⢢��W�N�Q+�b���q`8�}�p.����[" �(��f4L}��\�]��U���M"8 �w��m�֥�:^��k�F7�)�+m�ėo���Ti7K�*2A������~�#9996$�ٿ~��'�P[�s+��;1OS��ۃ[S���f�R���(�����| a���]p0��^�Sк��!���4�cM�Z��Kn����F�x�+�a_��IM������\�?#c��#++�_f�vE�����:���x��ZE��.��J�b��DSW	@영��w�Y�S�u��Dg��r2m��au��������Ss�l����͜��,�М|?��QSV��	G�e��[.��J�+ԓ����A��}1�Y25\�+VxS�07���a)\d\���Y"��.g,T�ݔ ͍�YY\D֙���ct����v��^��x
�,�#���xϱs�OO@����ۖ[��{�5�-;G�����E�i��G�#[�  ���y+�Ń[h ����6glE����z,��N�_%��������퇁>u���-z/3��sgEչ-FC|�eУ�U�顱��@KA��g{ٹHs�t���Q8��61t�6ko$�rZ�3� j\�g�V�Xa�$��@����w��t�w�UǊ�����Tˍ*� D ��}s�]w��r�G�F��Y$�*����0#w4XL���D��.�X_��3�j.��d�lE�{����f�O��hll����-pf�:��H.�fl5��8U�����,sG?N۠fɃ
�(�����ClGױ$�^x���؏-���;���f?��g-�OKJ�r���nm��H���i�[ڜ�vV��ꜱ�2B��F}0޾)����ǁ>I����|��r��ˋ��%N�ܥ��|����VP��1Jl���V2�-� #޵,M��օsk��$��1�)��r*],!������	ɳ��Ϝ9s�2hVF�D�ߑ~Pp��Xe�i��]�ez� ͓�^���xs���� ���pW󕖖�D�KNA�;������g¶���%^�&�?��M������w7E���\��  +ц>*b,"�#��\��Ãj�3�Y��c[.�b�b��?��������v�wĪJ�&K�j��F�'�$��TJf�6���c=��&�kO�.������#�<�Ӛ��������+��n�����.'��O\�������muDĈ���!�5�R q�D"�
}�[�`�~F:Hm��Q��T󶠧�Q�,����WF��c*J\�ۈRk�b��z� #�5��YjM�̃�ڞ������4����I�X7ť�$[l[qҞ����cb�*V��\UĔ/��u���RQ�'�eE�}�����˥�q�Ôp�l���&��G�V�ǲ�v��_|�˭��>5����ig�i��r���@A��6��	*N�k�+O��t��%5k�Pv:���"17..�m��H>��-,���M������9�?��/�병:���e�,�Q	]�I��k'*�,������"�1��/K��	+xLɄ�� �7����m�W��8���^�mm|���������x��P��q��� ]��|iU.���?3����=QNb��&U��H���6�J�Ӂ�3F���xxx;E&��bw�:o�#I��'�o/|�0}�/����NC`��nٛ�D����\�LǸ����'
�1[obTbq�;�{[���΍b����x!\ _�hl�tE�h��:��ٌ�<��P����7�gM�@�2�S�p�Umŉ�]$"�^��ޜ�����l@&+**�	vn�����饥�h6s��~}���?z"�b�4��2{12�7/�|������E�3�=ҳ���B��a�i���w,�(-��7�/����L�`�kz�{x��##KvZ���da鋬<<t�>���ަן��h�.-@�:�~*�ʺ�o}�D����*�rz�k�}{�y��S�*b�"��HU��I��W���I�*��K�p�ƀ	���n���_hg J�仨I�}*�#�����4ռض�m���⼴����
��ws�r��5��d2�� �۬�?�c�ҕ.��L�X�)I��&�:>^��&��}+j�vd�L����Alŭܖc=NWFO�#;��	 r�q+k�0�^E���2��G��񟐜�����X���l�;��κ�4������W�|��'����lB�#���.��1-wH�Mէo�˄<Ѐ�N��!`�W��NU�m���%�F/[&�BA���m��Qk Y�>�彄���HV���k��(+`��-��3"�������`K]P$��Ь����D�ؑ��10���iZ��j�">@L�&�J.�����C#��{����;��ڼ|�yP*���{����"�	��%�Xׇ�!�e��)���k����*���أm�~��������V��D��Ϭ�N5C��wv��3L1K�_��x�{UW��S�ȸg ������5�?��ɘ����#��\�z��-�I����=�@jA�����É%;L�������)UI1|K�����}�9C`�~&%(�0�.�
�ٚd�ܚ�)Y
T��~��0�"^a�>�XŜ��@�%�>Q"�J�B��DL��ԙF����|$���P�Z@���76������)��N��&��	n�Q~*��￙�j�����|�)�Չ^i����:3YenJ��twFv��8C������r�`���`#A�u��#��/��J6��A==!A�l�Cx-���\�i�[0� ֥�hv�j�'��x��ㅟj�>�9�rb#�&'���Kd���K�=��O%[�A�Е6�5V�͡&��Z4$�i�ո�l�ގ�+W��-\sDq�}�u�p�0��V	�co�Yvs��m��5�%ٸ���I��0r�D�?�����b�9���Y�� ��bccC�u�w�˷�������TF2��1m����B����ݐ��{4�ׅ��">�H��p��N{{{붡ܯa"�L%⬼��k�J,����~�1$����^Q���WӏQ?Oq��n1��'IڷI��o��v{ۧ>�h����鵒ޠ'��E+A�#}$���o�����߈����:}pC�}ˉKVە��9-�裴9�'}�1	>?l��V��H�YHٰ��1�S@`fo�}�pQ\|<�䀔�hl�TxE��;}x(;�B�O$��L�%�?6�P__Lʓvbz~���H��	��0�%�j�.���`��7��G���1�|�����"��$���)����1�b��������9�s	�o
�
��k��?�Eyy�!��J�|���ٟEl�r^����x�sd,�n�(ieeu��;s��yI�T�⦪��>�۾5q����j�$����_)�R��bMդ�>�\��;��9^N�Dz�2;�[�:~:��}�����&  ��|6j��{�5|��>�dlYq�4���_%�Oݕ�Bg�o��́�S`�<K�D�m̻O}����jxX_�36�.��o��q>1)�=yO�S{��4��I��SZ�*��)@)wJ�rfOn]�;�g������)ԁ�q<���@K�$~�O���?M���|D�0R>�!?5	��Q�%j����Zg��{��<�\�[P#jq�-amN���U���56�?%F5/}�( l�я=����D��	���`o{n_��0J�s�|熹�IZZZ��,J1'3�b"�������� Q��r��g�K�Q�~�RLO�TW��)K�z��&\��@o\����U9�|6�+�V����ݲ��d` ̊�(< w�D�W��t�G��]Z#
#���ЃT�w��_i����Q��Lz~<���J�=ҵP��'�����/_H� �]�7Tj���2V�S��L���s��a|Y�ֳ���VhL�uZ�B}���s����&{�#�^��D��`�5E��\����Tsyx�M�.I�|1�s��G�*R�ȸ�bWlm��������&�j�z���44\ש
�q���,@����ј���VsW3��V�ޭ&W/�X?5��0���,%&��(���w�h���)�M}S��|���;0�C룚��p���ٰ�����{����K�+�z6.g_	�HJ�N��)sL�0��~�8������=�O��i�,�?���988趷n���AxD���|����j�������ǎsչ�|�)$��B}{Y�dK����6'|�a��(��b���	j'�a�;U���ջL'z��M�yRP�+�l��Q���$�S��lu�vP��r?�G��#v(�},ܡ5�9��O�U��MA�
#Jg�b7��Q~I�`���IHe�TS^>�Į.����ܽ�c8����nc�@<��L��ڇ])�Yx֟ߴ��V�W�\s�+J�:b��vq`�d-���
�_{��rt,pK��jqq147Rq3k�ZS��$cAN|#���~�|C���#f��n��/����SE������VHI����/�2X�菝%{t�Z��L�1c���4�_��vF��i\�s�����E��Y�͐����
���\xډh/�$K�U���iERu���S�9�o�J����vNjy}Е���\��ܐ�"h��$�yuQ&����6�1w�j|���>�i���2L��7t����^2��5X��i�k���<]��E<��$^�,���Dj��o�d��?�Xt�����%������[�$�t�X^^�]�����:�{P���(�N��>��#j#��I����V��G�½��e�Bd3 N�=΋8�p�j��z��Q��iaa�;�ș�L��}?���4��T֯s��t'�A.�k��������҇��p�=D&'2�����Ya(��S��b=������F�7���o�KF�M {{^�	��)����y�t��g���{Wk�>.��@,<�l��Z �4��f�*X�&�P�9������4�C��z��\}�wNT�S��<L9N���
����ӡ�I��y�Ax��újb���.�E��J�}q��e3fek<+�{-#:��H{yq@����Vyћ���KK�A���`�6��',��� o��G�KXGlw\Y��4�7���yw����% ̎ﰀ���|MJ�}����\�H�؟Y����l���I��a�栺c��J¯^��g�|���h���L��p,�S�v{���q�ē7hA��
<lm�R�H��wa}�c�l�b��VAn^��+�}��Տ�qk�;��V��X�
`D����:���������BrVS#��;B�L�i�  �9(�:��Gl1����T������;(h�f�����	I
�u�����}�m�~~=؃t�:O��i��&��&�bkq�D����hԪ�˟�.�%�����8֪W�s��A��+T�K᥅�[���FY ��w�F�k቎C�o�IL��U ~"��S�D��wu����T�ء�^��1W@��#3�]$9�T��s�1F䇸���m���.��F���.\w��P�������1`�L��t��'��"k*m���pY�ć8�����U��0��6��=�;�]]]���$3��i)�����y�8��=vdh�q	��xI�cG�&/E�E@^������t���0;�r_1Ҧ�	�Q���ϟ/ǲ�&IL��oM�{
��L��u�7���:�+�[(���ZE��DE�W4�(��'�5�{w��}����`���:�A�`M�΢��>@U�W�G7��"�3�0|\�e	Px���gk6��5���`I+�2�~Ocg�M1+����EW���E �����ee��4���,�c�AAA��j�ƈ{��i�$O����|(�y�n�bbZz��B��Yk���{�e�w�������<ǓJK^�VK&�`�1�S�|{�Y2�Y�(�c��mV��4@p<?�֖�B�F%����cv_�!�iLP����W���$ɂ-|gML���J8T/N],�M�d7�975t��|W�<AqP�d�����,f{�n�Ch�=�W�_	�[#�^�����x��ڀ�;K&�І��胣mj�!qw����'~�dwc�7z�A��ބ��t?��	�M����@��T���y�M�����FZ����i,�����(�p �����
�`�C��'�_|(X-���uh,��Z'�?�ځ�L~t�W��o����P���)�qO��I+�(�ơ���֥�ܒ���~�����lУ�����V��+�ż�8����	2q�)�Ѣt.eQ��#gqq�y��Kz�Y�= �P�6�-��5�x��OPk�����R�>�?�X �ޚ3����*�I��h\ N��Y�������ej,UY��Ej̆�aް�?tZn��k�^����{~�Z�$�P	�'���}�f15`�j�ܯ6�!wI�,L����&ͭE@H��=B�g��3�w���[�ߏ\���I��M6
����{�H�}ë,��r
	�:�m����% �Vi�\��1m� 饤���"��1�r ��y��Y��QFzlll�VD1M��\?zT�K�������H���)���iʈ�(;h `�Pҋ���
ƹywd$Q����mO̗N�z�y�u��2�V�x��?�\��m�����װ�s��Idq��;�X�֩8+>0�u��uը��Y1����p�U���-��
�C�8��j*�j�<#��V.���_���A��i����p��~��LC��6 0O}Y��z�}*/	s�4���;�q��I�wj,�4�g7��#I[��~�4�p�c2U�������g:7hH���c��<��׭5J�:��܎�}�}k�B4�Z��N��CXX�=�8�0w=1��P:MP���Ly$Ǖ�_H�v�at��g3�|3B3}� 3nu�v����ş�n���c�����z�e�6|�E���:��q�i�������I�=�ܳ�M�?L�ݥ�4�nB����������ا�O�_4�M#כ_?���tni�I����LȄ^Y�����3s�	$�;�����̮���m9c�^}�+�����!��̏%!�`����c�@��iٷD_�k^c&l�������P�i����*`2{���!%Em���Ƿ�K��S��UO�?��^�";�����H��AB�ev� "Cw:���\���q��<�_hq���C<9o�oU�0�W/Mq���>�HϏ����B�8Xǲ๗���cθ��2���߷�Ӑ�8 ����;�.\�RVQ(r��y��-HpW#U=8�N��a�W͛�Rw,�_��NM��`��@.�����<�SK����7a���BW�l3bM]P� ��ʇ����H*�9:+��j�nma�������ќ#9�a#e���V!�HVh ��l�)��I�u�<3�h�欞��Z"�rGxz���zM��}��e�w��Ɏj��qq[����D�C�2�� CuO�Yw��=�;}�T�R��fT'M�7r0�ڍ"p��^+�O����܊�� ��ݐ1>�z=R �?�K�����(9��������~�=�� ���Z��Z58|)1ދ=�:֝�N3�y��D9B�h���K�6t��ebT�?Mw,�l��JH?ށJV�q�^g_¾
_�QW%ïW9A_�=��9���Gr��⏜ZB�q���9�)�t�q�F���:�z��]d�� _f<���xd�L���>9��a�Dg�u����9��CVV���
v���i��X���SfC��U��a�q��Q��vp'q{�\�%����`�Զkm�`�����V������,bGY+?�-Z)3�3�^�(�
To}�W���No�x-=�x! ����|P̓ӄ�H̍n����;�`����:R��9��=e՗�o��q2�܅��𧱛e�	:J{���+�Q�z�i�)G���!���Tx���v8h$;����_�ulz#m���`|v�M�B�v�d�_��w��f3�P>ii[�1�M��'���.<R,�����;8���H%�v��<���Je&��1;��Q0r@��eH��T�sZ�-0��s
��v�r�fOʾ'��C#�ʭ�Gj�$�(s@u�~KZi.��e܅�^!�f�,�W)fV�c�V���:\�a�	A�+j��G}/0��m���x���u�,���`��J�4����c�������=m���
سV�S����=�\N(M~Rom�4Ec{h �`��x��"�6�Ǥ��	v����z0O�Ȇ>xꑦ`�
wb����]�A�w"�}q���[����f:�O�o/��3>�;'G�<�ä��z�T��5��h��L���I���e�e��>�����}�����di����2�w~��/ѰA6��~�����]�!S� �������&�q��ٓ��	B5�_[[�c��N�DPa�)Mǳ�v�Q&���D�_Fp��i��$SRR)��b�yz4�J��J�(��@�f�*C���D��6w�;\{{�Q�zV���(pG!x�d��E��o�4m����>�}B�1�=<16�.�Df���#&���vRVd��h?��b{��Q*��n����C����¡��������[��N˝a�h�T6��/"5���5
�geE
������ж���~~���&*J��~W+�Ϳ��$��KѰJ�l�����9��$��ZwBr��<�����HZ�s0�G$ �p9��#"�?��� ���&+��Hl�c��G��b
±��b��Ɛ������� k�4t�����Sw�i|G�um�W-15�S��G��Bܜ
Ǵ���	�j�X���,�r��j���� �*�@���jCi���n@uo�v��"���~\	�ng߶���B�ڈs-`U��oa�18?9�܏9�W���̱�;� o����[���n�B�nV]MM����^��l�����klJ��i���3�h7��n��3��Ʒ"#��r�2еUw���z��Sl���}�'�(�<�d�j��3�{NV�p�hhdȳx=���>��zr�R������VHM&`ݣ�N�Ed�?� ��&ѥf��2,7���]U������b��	���T�%�]̷_ɕ�;�?-C6�f����u��WV�9���؜�1�{7Xk�*>,�~Q���$aq�j�\�Z���:��s��)�����X~ԯD)�k�	�-V �r�T{�4t��C��%H@X8�M������"~Qz�'C�����S�I��e��|�=�_��޶NCy�FA�b�r˗>O�e��,z�D?Eף��'L�6��C����ق��$OҐ�!V���m.��@w�G�~���B�C\��C�#,�@�LPZ����0�v�T���R�P�PճR숵�raf���{�5�e�m�u���,��`x�]�P�A�i��E5��4,ߟ	(Wq�J/=��~4m]�U.J�1�+���g.�.���**M0Z�u>�s�$՜{���v��Q|�S#��پ$L�V��"��*�q��4�c^(��~' �N��#��8�*`
���<6�|���p��n�+��7`v�>4���0����Ό��d2��lÜ1�y3{��Wc ���O����JG7��/���ן֝�BbG��a-/ŝ>��gl8��'u�N	4����~��YGYA���WQ	���H�����'��?�C�9���M�ָ+����r�,Y�n��'s�,c���;���Ii����P�R��������$/��N�>��Þ��h��b�\Jܸ>�l�?S���(hl{U�qR:$���ׄ�����/ߟ��]~.�o�u�Y��"�#m4��ۿ�JJ[�nG�;���^�HC��u��~E���?�?2��,G�$i��bnͳ²31���s1]��<��hV'Ʃٴ�1�l͙bH�;j��t���B�m�_���Z�q�O��1�����;׌9!I���Z�"%4��M�Q���m.K��>?UvJkm����9�#v�agc��[�IWCC�k[�޳z���[>���1#��xƥ�Z�2w��J�kb�Vv;����.��rxD�l��`��ዚ1�\�3OA�ZZZ���<�I�=�Ex6;%� ��娞�h�8[��+��%�
�����;s;��|n>Y�� *�VMu֚��p��8ދ_�I�7�!{ qw0���SڥN_s�I��;�����阎��w��i��g.*"ۮ����]ŏ��Ȭ,Y˺�]rv�AlU��������w	�o�d��׉*:��bM��ݡ��k<�A��U���e�j,�z�t�3M&�����Z���ߋT�N�ɲ�b��W$�RW�%?��ԼH@���|�A�Gh���py���������D
��]"˫�ulZr+���H�s�T��1�ϥ8OrM�7��%�'�5:���^�R�!�@�����{f��2�����£b��Q�2�ؙ$ҽx���g��)^�ڷ�oy-���+����Í��}�ظ��2����$9yx�cBk�p<=����m2�zp��Q4�
��}�ݲ}�Mv��o��$��;H�޺����i�W��S�����T��_���ꣁĝ���`yi�f��cONs�����Q��snL/����ͫǟ<�Os� r i���훂�������4j�e;�U���tл���ɋ�#h.�Nc���:��"�axdda]��:���n���4�uZ�V��8�"o���$4�䓡���r��KI�x��_|�{��8�aw͔S�%u����S@��@yh��a�}�?��܆�z�F������;g�8�;�b�5�� ��psn<���Yr4;�U
ܑ���g{��Wq�֨�����)_|Gl9j�FǷ�K�+�]~�|[�L��p�ߴ��ڲ(�������}��.���ut؟z�!�I��-A�	�9ո\�碣]���Y[snyYJ�<����W�a;�*��\�@/��Ų$����yO��@�O��hh��Ԍ.�<x�=���@����I�Ʌ�P��4�i����/�?�; �of/�~����³���xGkg<<#b���caa![�bE�˫�vw�hM�Լ�s���ҡ����-���R�q�C��1�3k2��@,��� ڪ�2s�=L�5�\������s��(�D�	��n��W��]��n�r#E�M}���7��ݢgԌ��:��
E)�����ɦ@���j�������Uꂀ�*,q����2S|�>y1,��Z��S�F�S"�c�4?t�\(����s�%|�S���o��e�9{Ѽ� �^�y���˧��n$(/m.�As�S}Hb~�}iq�,u��������V6Z��ܳ�k�xf�mK��aWeh�����wu�wR�If��P�Y�Y����0h\����Qw�$*���)ҰA�]c�0��%��"#��F�k�8?8%�����3�����d=����j$ԔʥRO_?A\Bb`` �Er������f&_)�L!�=��hydYHn���~�M����L�ؠ,�H%����t`�?Xb�Uu��� �ao���*��;`K�!҅�g�2��'s�sVK�r�dC[�!���V� ں�V�Z�K�H]VV����2n�K�ݵi�H|G���4[�ᶻ���oc#���>52�51GOE�kfh���2G����޿�l^u�6�ר�����I���Z��ighJ輻�5�M�;���:�Ö�g�C�vt���GJ�l�� NN�(�<��+Iv;[oΏT`������ʢ�Q5����؞d�[-9.6�\�Q���Zφ�<��������}A�����=�B?R
V]��5 � � ._U��fݧ?v�)�뀫�bԝ�216�y��A�5��ţU*$n�gn�`�����իW��� �L�R]s������4��S������^�e�z��PC���?��x��Ĭ�W�����@֧t��d��������!]	7ln�`>{vhE&r����\�c��'��8�"���xp����&$FF���K��=Е���lii�T�*��H1z��D"ָ��F�:�QW����iȹ��GETz$�X.t�l�Տ�;>�g��+��{[�m��2��A�ZZ1}G@�e���YL�p\�* �H����׿U�1��\�^���*��׏*ZV+k��/^�---}�"`���kL�4[:M��QƝ7}�����َx5����<'R���r$'���Gs����L���Օ���L�S�!S���v�_�C����ٽ���k��me����6NN�GGGׯ����y{{;���;���$��±�[�� ��a#���J��o�Xo@��Wz��**7�o��~*(,tݏL阅���>5�,f��#!���߱(��\6�"��J�3נ֦�;�X���Q.������hGG'''�S|�#"�/��P�-��h����j�c�S#��6'I��"���Յ��KE�Y��E�#]���3ϻ\u蛡� ��F���G�����������9����@��N{�Lm#���5O�_M���ڊ���o�z+��y|�<e���G,,����n\��zf������T{�6��� �o�����j��*oP�f��N�3��LÚlG'p=11���1�=��W�͙�4�a��Q.���_����P0z�{O�'f\_����
��:���\aG��K�+V6�8/�����;/}��S��N�ٙ��?X{�e���,t�g�{��"�M3 +�TT3w�S�B��-K4�@��Tn���o.�Z��	 Y]��,�I�טE\�������w�xoWd�5���s���㯞�����7Z��"�>��jGˠ~�u0Ah�k�<|�^.T}&�99O���틞���bb+c����G7�O�%^I������@A?
�/����L���7�$Q�GhM�Bگ9F�]��PhVͻ}��i
���m���1;~�������6�c����:N�=�Ј��� *
J�����}o�EU���JǉTp&��ǘ�0X#<)�}�d D:�x~��u��	 ������T[ϼ������6�BXR�;N�${�ul5�2����<���Y5Z�����Lb߉%�9ɩ�I�n7k�j����sI�+����'}�BDi�q����� �z���aRBZJD�D@Z��F)�Mw���l����DE@$6!nR�- �����|��k�sTp3�ֽ�{�̚ƽΩ6���
Q���v������Y`4������`�}h8�vw˵���y�b�����!�A��d�d�IQΝ�w�W��<�QG�rEp-ź�eIA�w�����Q���%��-����E��v2��;)��@h����/��%jY6Z�X�SW����Z��#GI���	��k��Q�v�9j��z���w�T?�W���qE٧�W�VW�n�@�F��<�)�(EI.b�S��f�A���k%[�"T����u��	������C�\�5�P��,!
�$����ö�|&���R�>��m�E�+�&S�ʕ��ҷۘ�	�2�<�dx��gp�R��oVW_�a(�a�䗾>6^��y��D!|�!�]��iC�'��f�5U
�6X��좏����Rj�q3s�����;Wάx�%Oj�2x�S�M6��������K1ҟ�73�j� �[�'�����tM�"*TZv�K� �m 8���\R����5j�(r���A.��MjР�eM_w�v�*y�p�\��"c���M�5�����g��+,++S�=�O�S�1��T��d��]Ac9Ӏ)d99�_>݋ �d��$�0GX|J�%��f�kuI�R���s��op�ۼ�6�֝�1��Kb��갦553����˪�U+���ګ];��hZA�����^(K ��r���E���2����X�^k�}��WcQ;�)w=�P�:��J�!�u�3�fNR��.�vnߍ��}Ĩ��#^��=����Էc.�!��X���)�و�n����u��+vŬ�hڝ�R3$��G��Yӥ��6�����Ư�����g��v��8͊��Zo?�a��*D
�B�+�*T�z�EĲc;�R^n?U�`͔�h��@�kG�$q�ɓ��N ��K�@��Y��<��@��ڐ��-�I�a�r����s�s"��[�a��Z���;�T����+���gR˭,F9�w��x�~r˃Y�t�pB���l����~�:��p��/K���*�=G�vM���D�][L���r@tf��y��%I1R����`!�7���֗0o������T J�{v� dle '��kl\.O�k�E5[�t ��ۨ�ˉ��z��>(�>���ш�����������&�TT���*��Z[���d5??�$��t�p!��epӊ:�/�ֱCb���[���[ќ������r����Yf��g�~'��ss��*O  -�0�:+�<��Z��^�oOOr|���z��;0%�m�����|��T���ד�/���d`�`�|gyhUQ��AHD�
����{_X��<����|��M�i��Hz1@0'���I��~���-6����0(�:����ݲf�1��'`�x_�3�%#��D 3%����ˬaي�~�i���F@m%ɎC�;R���p^�Z�!@{g�)Lbq��)�J����c�R "�s�V��C��0Ϫ�m	b�/�@�@�@�Y��n@P5�.��cT� l'�>�4�k��'�W]�v�(���C�uT�j���h�ܱ���ぐ���S�����!�:W��������Ӡۻ�V	;��I?;����5��~q�J��"S��~󴰑�A����P�~E�����o4P| ��=��m�N�ΐ�q��=8�V�S��k��ؿ�зl���v*�j5n�#T�ǩBW��Řg�Vpp`m{���k�'��ME�}��.�|��|�w؍Ilu�s�䭏x�#o���:�]�_��'l,�
�M#cɺ�+mv��+2&FA�0���v�jh�@�14�]������U��"�ⅆ�0�q�<�oS����|��cg��B����	D���w�/�aW��������
�#��-�aZ��45����O88y?��8wnj@�q�؛�" �{V�{^�N���n�~�`�<���^N]kkk��N!���x����}��R��<<t�g�����jqlJJr���о�Z�x+2���n���eIq�
D�� E�c�3NM��fWW��;v|l� �Kߦ����u�(�nX˖�o���CJ�R�XY�2�N�o<|����Ttё 3�����@3��� �c�UH��|�MI�#Tc�-�f��#w������1�NV������I����s�Ͷ�U��ᇏ��Yy7(�M̩?��a�*�3�I��O~S-dz˨���J�)WK����
T��}�"�����A��s9jק��4�vIC@�ʁ�SZ\���L׮Q��H��j́����+4��g~˼�\�m�1�Vju50c���93��EP)'o''7>���J�2@Aن�[� JE��~�s�����ݫA�8�o9>:��=]�o�+��l?]��10� ��* P'�ù�Ӑ�W��ȍd���k�8~��P��Ic�����r��G���}[Z�b/��P
�� 9��;9i~^�N�Z�Ĉ��������>Hao����	��ۃ�Ji��Y2	=XW�wþV��q�L|)kS�L~�����9M���pWS�܃:���.��+� ��n��$�8���$�5�`������څ����Jok�
���'8g�w:T�?�Π˝�%j���4���N���F%�:a���ܬ���[^�n8|0O//��(����:(��5N2���3@h�H�;�*����:���a[��s0��Q�GÄ%OφF��g�J����? ����kV��K,��Y � l��	,�o���a816ZqѴ����v���)t�*
ID�hX��j�S�AK݃r���b���n�A���1�+����7@�4����yH�<X{���z���0�g����'rr�P�H������P���vv��߂ ��?_�Fz}��ȻH(3�'�d dñ1m����x��*���Y@�Ђfn�s��ppk�� Q�5�s�����KK�lɴ��׋*U��28S��D��%A��#���~�f�?~���w� ށ������!A��=T�
0�
��8��۞_�/�<7%:��IgC���6�Ɋ�'�x�2^T=ym>��r<::z۴�b���g�e���貇h�j�P����g��KH� ��RU�x��q� ~Z����M�c�
cۜ�+�υp�Gt���6>1V�j}��.}�]=a�I����Uo+���P���qPa :��1+&�~~���PJz��]]ݹ�O3ϑ���箇V��:�����w�! �K>��m^�JVRb1��llo7Yt���6��#�2X;>2���N�|���v�3�Q�[ݴ��Ő��k������H�B=�5eF{cZ�7f~'�b���Vg�^��[��)�/�{��[�'�m7^�[
�JP��<�Df���4j�lt��Ҿ�N�jg��D=�5��>���?��8�bX
X��_����C��b}������ �$k9����l�� W�B��j|_��)~��Q�����Y�ÄG��o�]��-Sa{���&�}X!־��KÕ�vxv�1�3�ԭCo�Q�[Q����Q�L���֏&TM��eٹr#�)0�~�~S����TV��2t��
�h�n�SqB���\TTJ� ���-Jj՜��.����-�C�4�7��D����"K�(����ר7n���X��-�OІm�����@�\\�A�����ly���� M��p��yoooh#U��)�lm(@�
.���t�
���
C�(��2��RΘ��Es�0H:׳��R����03\�]��Ó?>T����: ����3#ğHB�����G����-�k��TkkZ.㣐�AK�W1� ������oCű�'�9;�>&p���:70Ѽ�ϵ��l�u�B7t��I����ڟGx��p�J�:��%x����7��d|�	@�;ЫЎ@�I�K���EfV���I��;a����k�*����. ��������&�(���.w����*� n�pvgk��4G���wS�n��Uᜉ���241Q11�=�
�a,t��p�������&��H�AT�SκIL�]b�c��O2�s.��������H�4�{p��w_�������=?1997��' ��i?�4W���o��Z�%�H��#�?`�jy�<��+P����JaL
��[��*���ӵ��S��Nש���3_�?z��a'��������Rr}����tvwM��mhh�Ʉkk�������yM�1.�L��ӆ.��w�D���R�؍�+�m����%���'P ��6<C�끉}W���з�"��@SS3:]�w͖V�F ����!�XP?��j*��9�΍�c~L>�����m޺�3��ʻ��Z�9�o���_&�-�6+)+O��'���744uudffg8%l@����Q��ķ�6:���WD�\��ep�����6��P�V��R�3T߭��X���y����:Z���a)����5fL���0����8�&�^%̂��
m�9$>��cs?R{�s��V��ON;�����)��@��zQ���)����iv�Pi�2���c���ITT�9��옘�����������c�������l|z?Խ�qYRH���= 2�m�x:1 V�o�PC��$h����u���Z�� E�d�_������񝝽׸��'^�m`�:i��u���h~�t�C�L�?���։?��i�-�~�+�(�~E�JY1��VO���t)��/m׷�&��P`�ꉵ�@��_.�F��r� �.}ئ��o�%�@��@�yk�N:�k��]y�C��������k��0dB|k�6e&��~7sM�����N9 �|9�q�2��ep�ˤl�����w��b?�5.�S�*@\���_�hR3�T�����[L7?������r�pw��D|�����S6?1Qt?pCy���M��|�I��X�f*p3��o���'���1����.p������]��	�'u�ܱ�����3�Y_o��Hl��c9�Ċ��|q�A:��Ί��]���c�{�`rS�P�SMr��ȋ��,ǋ�Ϡ�H�V�!�U �omm������p����:A/���d�y���Q�F6o��`*���ｑ�(�X���dn���������9�}Z�,P`Q��
�� �;��7F�������B<ζ��SRRn�(�������c��%;���ڀ��Vș��Y���6�p��oRp�>Z�@D/���a�kV�frV�;w8ZעWƠ���<f��y��cb�=6��W}Q�M?,8�h�HB�$u:6��3��_x�*���ԤT�6��9��A0���]*�`�T��h�����@�3�r�@�ж(\�f�̪]�!N�bv?�I4���5_���=����v�T�.-��s��1����9?T:
�Wl���5D��k�^Cc#�U���Ufqfff=��fM?�Rg���#�~��lvՎ��՟���t+/��:��G|�o�[���!b'k9}�=�eU=c��j��Jq�c�X������OLOg
552�1�����=$*���K�$���Q�K���)޴�՘/I��sT/:UNUxz$�?�377E�B7��VsTVX��l�jG�������g���sq����[[Em3�sB����:&��7���Q�9�C�@C�p�j9:>V�C����}��h�X`Qf��c����<��Q������ă���\'�4&���������x���ٽ�1��h6�w�ޔ��g~�����߳VU���7w
E\�5اlnn�O��h���@Y�C�Tyi�F<��}�ZY999�l�G���O"��%�+�F�摥cG���T��J~��YBozf<��Ϙ�y���3�qkL��烦��خ������2l��oSxW�f��������LYV����V�%C{���s��s-E{���A+햷�8��s���S�U��3��������+����%�
�''g�R���үb�%���:�f���W#��[NMƃi��z^�8�M�CM����S}��FyAΞ�9�@�|ms`9�ҿ�-8V�^t���Zƽ��Z�K�΀�9Ѐ]9�I���'}+�g֙ŀ���+�f��|_q���*ooG�Z	�..."��\�d��%�3�{�z\-���yҜIݰ��6��$��g�G]���iT� >�n��5����� �yG�I�߿�<�Q��q��z~

=����i�j����7����Zo 9��L��n�_�o?�ӥ
e�Q�?�z0I�G�/��������eGkk+�i�Q�ؒ�їC�[�}K{�4 ,��/�ЦU.H��^gr�{���c�����=�M�T9M�3�ͤf���t����M�7\��j�}5�����a�䰵�uYU�V��
=M�T^~b*�b�6z���/W�gA�y�;��`�'��4z���i��Fa�D����z����˹
��1C������,-����Jf�(��"- )7Vc�����[;�g�g����:�lub!ߣV$ظ�0�z�{��-��&�9'���ΒQ24J�yZt�>��12���;cE���2F�V� @n��Y=	�|($TVS�yu��ЕE�[��ϙ򦁥�:(S[[[�_H�ek[��@��\(&���[��@�Kl凜]wou��!��i�<��w��\vB6B�xn@'��HB����^������b���aV�Uz{�C(�\9���KU��
��+���u��j�|0+�.q/���B�k9�����:݉�!��ϼ��Fr���@���wa���u�a�m~vw���
:ϵc���F<{_P CAA��� �z�8�)h`J�uZ����p2@���u�+ukM[��<�6V���UX��=�J�?�<�)�M�ϟ��@�&����r|���Q�K>�-�i\�B.�"����$�=�	�^~��Dl���,^,�Ie���}��f�|�V\�	�c0��گi���ܦϋ��KoԸ�;�~�Gi^��~�|��Xс;�8 ���Q��� I�Ф9�^>֘���>h��P��ܝ�����F��U�p4��cL���Qٯ_�b�KU�7(����By�:�T2�s�p蛜�w�?����Er=�)3@oAiv�w��D�c@�{n����������x0j�eH�4@��ԋ�ܜYx��묟�ƫ�R�F=c��;D���r	��t6���j-;�q����oҢ����4ϣ�a��U�۹�cS�`Ri�ݗ���� �)|�R��~-W�n�5����(��峺�v���s�%k�"#cc��k\B�l��s.�l�c�8Y��u*�P��.~69�[�U�~S����9�V�d)iiPf ��;*��l�A�//%��-�	��ß���T6�A5K%v���6P����A���ZU焻R.���`�w��^��1��!%�c:9��C�	���CE�T\��rA��ކ�5%�Q2�������vߣ8�?X�`t��*��~���dT|��s���
�CpnJ�bod����z�D���4��$BMB�
�O��S�UM��ߺ��Dn��p�z���籢~pj���K^�NqT��z�	)ݲ�����.z�Ey�辜4˕�k�x�5a����5zU1�$�=<t������XR�L ����̲6ϊ����蟼?G&�WK@IFūA���b�&��F��*��\�m~��~��xQ��-w�o ����ٿ��V���v}Lļ~�w��v;kț����o�:Ď��e�5��@B�7"Q/�h�J3�["�Y��M.��_L�ݮ*u��@6{hp��Td��_�D�Ȕ�ۇ=�������⟘ӟ�*�\"l���J4��a>�ք��mU��G[HaM�j	*�ѽ��_�����34�̪�ǰY��Vm]gb�tk�6� 5��?�_�]�'��^���d-����T���L1wO��Re�.�T�p�K��Wm�;���~��GNp�f2I�����v�t����ᗁ�v���~u������ÒH�ƃ'DE�ָ�%�P]�j��0L�1��~��D7�J�4�y}^rU�wf�}跲�c������˷���z1��\Ͱ=��	�A���BϫV�]F���e�}��m2���-���kcb�V�%���0��3�(�m�4������i��#yM�Pz�������԰0����kվ�*=�j�P���sv98�#�<��O)mW�w]v�G��5��=�\�7�%����<;ޙ�@�4x���C�c��� ڵJ�{KC3����38�B5�rļ9�v�Mf���I�f@Z��k����*��8*��d������1��r*5��0tJ"pbzU�8##��㳛�ț}|��e�w>���@y�?]��/J��Vx~������[[�|�〭A�^��`-/�l�}?�>�@����4��J�߉a�7�#W�ԃ� d�*�V���P�by�~ˈ��~��[%����ܐ�7�z�aA;݌�Ig�W��j��6�ʰ�Ȍf���Ub�gvB)��,]��-h{{n^�!m�ʔ���6����������+��&�K��m��J���K���3��_� �֐���qj�l��9�߈�J��S�����Br��V\����@����i�o	R�����1�{h@�C���������V���gn�E��ۋ�r��_�SǾҸ8���,\�A�}a�W�ȴ����u$йPa49��;�w�)P[�j�4V�;��=�vC�83�d�X$�t��4�m� ���''�

*���JUq�����7�;�����E���n(��n+&I�#0۩~�����>G?�VH�qO����>�
1�?�ׁ�K�R�iv<|"��4�ka"�8��z1&6Q�(EI� K\h(�
�O�GԒ�V�t���K�wrw��z�TIݶ7�ᨋJ��O��Nl�yLOm���w@�x|b��r p�&Wb��4A��0���q�ʕ6�2X�����t���@jL@Hkjj����V3����ѱ�O&�.�(�Ǯ"f��t%"�ľӊZ	�?'�b=�3����+�3G!ۼ�ڭ�Ɏ�S�c���1m�Pxm��cgg�5Lw}%~
���}f��Ѧ�;����iU[�Y���v����?A`p����C��;8L��U0��ƮC�rzz魭-xU�_��}9�o� ����2u �B���h�k�x�����`�D�//�5G�{���bR�XG�)��i��p�f� ��F�����*w2_��ZUg�8�Z��� owv�~]s�����G�EZP
�����&D_	���϶^��R�;���?A��7�|_��Q��<����Q���W�cp˻}��w�Ӛ���@R\#������ ��C��(��zc�||v�z��C��R���7�T��z�1_C��^����7wϯe��3N���[��w5Zι��Ҋ�A6���(��<����{�H
�&�7��:��O�/XR��� ���ŋ��A��&Y��?�҂<�7ea�>jr�i.�� T.b���O��q���y���4#$$,���pa� ������<)��ќ�o�m˞�6d�ui����R�xM�~�@+���%��"���t�>�V�/�lŗ���Lڶ���n���]�R�y�g;kj;n:�E�c�Ꮵ;O�Sé*��ٕ�|��k��t2n�sH��Y�W�tݔCf����.ccTž8�#%
���u����x�k�μ���Ey�O�_w��կ�Pl��;J"x���[(��6ǳ���?�r7���'g����ߘ��m�93���L�-;�؆�ӧOߨ�zušZ���)_��bzܝ�r("	c�-�#�W���sg{��^9�Zv��-RRRBF5��XkC#�����j9�����F�P*1[*���bS_��0�ޠ@�m����L��fr ljjj��g��uj��&�������c��lpn������_Q܃g��Ni�d�T���j}֓sC� ������k��S=O{��"O��P�msZ-�H;��n�1o�)o�I�53^ll,C�
#9>���e&�RY�gƲ��{7%ɲ�PK:��t�J)���uT+�h�OM���AC��U�~��m�������kW��֖_@ ��/��#�O�/E�\E���:&H(��\��>I,��UQ���Y��Ls(�=��J�R�������i�\�M�Y�~��e���A��~�t�6�!%�L鎂��vz��g�m�u��mCرv��T�`��2m��`�5۾�+��1P0�1��� ~O�f�C�+�*�H����V�n5+"�a�e��F�+z��]�ӹ0�X�Q˾�@`wA��n�Tc�͉�!��-�ҕz� aI�\O�������Q��ks�\$�T����b�<=��ʺ���~r�/Mŝ�bV̉��n�ڢ�ĳ��Ӷ�y�ć���?-�Ҿ���W�.p'|�{�;xCt"�$L��r�<ԋ�~��\��N�~��hy]�g��A}���o�����a�s�3�n%2b4x���7Zg�665�ttZ���O�#}���(���/��R�f�!h�~t[^g=B��d�'��_ؾ�L*�}>Y����0~�┑9���X�YE*�KO���-�_��UFK���������pS�"����204�98��Y1i��q�vh��Ko2%�<��=�An=�� 1�˖�i��f���0l"C��]F��:�g���9�К�>{�7�$~�	cA!i�e�<iT�i0�p�!�I�pO�Q��x%�'�2k���զ��$�R�YxVz�����
BV2O^��PS��Y4Mp�T��7�q�{�,�od��fTIiT9�$�-م�A�v�mUeˋ,��^��`ꏞ�����.{�`NF%������y���z��o�1]��#��"����9IhB�»S�S
�I>�%�u��A+���9��f���2O^��˻ h0��V�nX<�D���o�
�Ka^�ċ1����>I�{WX)�ݬ=�]���^z��O�w��}���q��!o�fƵ���b�"�τ!��ymy�-���� >�*�W�X9r��e�����\E�i�\-)�_|����>������=�5����ig2�z/���:�1��+O~la57E{�JT�]�sX�/ ������:�>W�vW����Mے��
�`V�<'.��������Kw�����m��&��xF��2��J�zJ���]N���N-@��0�����|?���#ؗ.ELp��;O5e5�[�Z.���".:�I�
��:<=�{G��:��p7#��`>[צ�X�_h<��˲k;��RG�x&.pA�]�U䎽�Ӫ�������c_'����M뼊dV�s(ܼ���(��f�a�>�Jmd�Ã�!}��m&�t�	�ӷO���e��'�uu'���,��������f�b�_T]'�A���@��l���I]N��x�y�'���
gN�u�����wI[^^�o杻���ΐ��v�>��j�VY㘭���=��c�Yu��nAU��C��.Ů-��[�n���K3��Z���0d���E���M�>�/��T�ݐ+�#���DKg=)��ʱ���00���ĥ!��km��8�m��=�B���^h��=�}������)�ﺦ��e>��M�T�4��x�H�_X���#�=1|����?yZ���H˂9ʲ��.*b���z�H[[[��
��0A����0Ѹ���>�ّFˢM�u�n�F6�����w
��,F� q�ɻӁ�C~���13c�,b[!{�|
���~�]���Җ������)ACG�zZ������o���b�Aھ�uӲ��҅��=QQ�M\���G2_�hlo#7|%v�]Ò'�{f���Zt�I��L�����p/DW�V��E٠���ǟi,[`�;��<�i�#ɚÝtg�����i��b�O'��6C�����Vr�ӣj�-�H����R��Y[c� ��:������J���������Ғ܏�_S�Y/ϖn����V�)fWZkpg�������ݶŶ���  ����<q	}_s����
�tɨV���)J�'��|�{�9Ue�(	.���8G�d �)f�?��� هl�v����{r�`�Y쮖K�x!��H���Q<p����%���ka��)������;-��C��M�^t�|�� ��G3��aJ�&��b��H��j����p���3nv�7���$��г}�l�5or(��6��_`X"�B=ww�ellL}�v��23���Y����c��O+�i�@z^�}�ЫĿE����-ڀ?=8/i��nɼ5�tww�g�.�$t���cCKC�� P�"�R�9�Q�G[��I�^�z�Sqzyq�H�ENqߔ��(�Θ�Z�V*����(�\�ş$U��-!k�����ڑ�d����7�.*����X)��+�4̜�j/Q�
� ��ҏ�Ҳ$?�ׇ�0;5��M�ԛ�`��'���V�R�-љGeT�+[p{BlU}Rчe��m��n|�H^��J��O}S^�(��O�\vZ�����I��r#�֣p��i�6��ٿ�C��?qJ7)�{X���y��}�����*�=˕��n�w��H�84ivA��x_�d�=�rH�g�4���j�!4iqþ|�/$$t4��Ԧw�I�݂w�6��D=N�Wf�?9q�����x�/��5��2~ϓ"VE��󇎎j&Z���������j
�6ۻ���.q.LFd�2a��Z|���_��
p,�Q�Rt{�Z��w���{r<cn̸~&gܼ�[�Ўݏ���S۶w��%?z�	J��[_�q�_��d�h[c\T�y�q�`a�T���)
��!�x81e����B�|>��an��#�-�#�z���pU�ez=Fا_�m�ުZCwAw���r|�Iد yȑ6[I|��c�>ߎ��}G���n�3j��zOOE�J�Y���J�U=/�4���A��|�b����>%=n�������RVVnv[��2����d�.Ցʒk1Y�R���3�#��(�^z	1x���,a�J��x7v@v���$�.�2��}��M ؅��
EZ@sI�O�1nZ{o'�ƿZu�n�E��@B/��mX4�E���X���c���ؤ�� yY΀#i�,'����4��|�$�Ik��1b2BsW�HR�
4�5��Y��a����٦�5�"	�}/�H>fA?�H^�\��l;tz���?�6�u8�������p�gMz̚ԣ|�#��v�-���{b������������~p4��yUj�{�^��x��;9;���9�
�H3����ē������Y ���O��>y��	:R�����tz��YͰR5��K__�
k�ͨ��E���~�V�]�	ь_p���,�LT�@�t�m�B�*n�I��0���-Mw�88��q���Q�V���Q�^7���<��Jw��v�������P�?}ɋ�in�e� Ģ�"�05�U+�۟�����=�� �FC[h�MMM�P_�%��=�H�t�P����`t=6km#y9�@��o
צf��T4�KWQ]��ӐU-� ����b%j��B¹��[�Ehq�bTX1���� t���sIO�kҝ�.��� Q�OJ*|�	/N��v��M#���bE@P��j���i�Ċ��{�z��M-6J���Ñ�8���F+3���i9�ݺBL���������M%�o��%`��wc�}6:n�����e�Fm�`G��0�e��ý=�_�>%����Ҟy�R�~����$�Y���ݾ�5hn��m?���q<ck?[����������9
0�e���cwZ�p������X��1/]�>�$CL�8���w�4��K���3�ݕ����S���2�����#Tsgc;F�N�-MP*=�R���S�hr�ѫ?B���ho�5h���Y�1ߵ�ӥE�'Ѝ�h}�[?e���#�@K<�H��S�.����g��~�w�l�4H�[	Dd����ѝ�x�qy�JF	������4���w�f��o"��4��J��v-�5w|��mN� �� ������{Z8z�̽�a�������E����R� }��=�qooO���N܍��»��l��K	RDh r���Ax����-.jݩu��_�Z�fIF��w\�u�+9ő�4�wo��D�����T��]K����F�+־���4r$���T����L�f�z��~�bbܦ�] ����p���qC�ZbACMU3�(��Qc������F�%�i�i��~�◔�`���ˋ�0ͳ����Y������;��A{��kǙ�;˧��`����E)�jA�J���,wq�j�k��t7p�3��)RA���V���'E���6	�g;]	�KPa#�	������*+m��#R͝�F��U.HU�2a���F ��47�G߈ ���;y���Vm�woe�m��4ޏFS0"���~�ES�<¶jSS�k��Ѯ«��)������9(2���$��`i��}'_q���M����"wp���ʟ���hoTX�����|��J_������l[���~������ ��M�Շ��P�|���B�C?:�ٟ��V��/9eq>.�-���ͤ@F�+��wz�:�P�����9�y.�L�S�]>��0u/:�o���R��� �p&̞��.�r͕�a��l���u�)<ok�G�Q|��]ϙTzQ8�w�=_D�A����.c�呋�P����a��t��y�Yr�L�q��L���/_nX>����3���L�0ē��4��*K/��:55F�� ����m�Y3�.��&�;&D�|��������s��',ͱ�5!���j������������^]~c?�/j=Ԫ����^o0uR�Ļq��5?��J3�p���\���~Xo�l���M�R��Dl�GX��#��q�܉�g)��pzG

5
�jy�v��a�3
�5r$���i���vO���H��b�JF�e�>�����X��~��ٶ�}K��4��c�9���CԔ����wQ�)@#66� �<�MJJҘh�Im6G8>��Z�Am|{�*1��6+9ײ���F�^��ZMK�u 
����=�S����~�;	]�G���﯑��Aሔ.��*vr� ���@���<a��0�(����~>?w�k��'%�?*Xͪ>}��gAp��޷��#8n�h��z�$�/�5��������S��۲�L�#dI���.e�p{^Ua)���y��#��4;x���㛃>�]�m�?��@���*����O�11�7A��k٨�&���YZZ���ׯ�@����;���5w���5��VcdO���Nf=o�4������p��7�/��7�m��Ode��UF�(a�h�=�2a�~�<p[���r�|�*�������.�]O�t��Ԯ#�q��rȤ�0��0�Q��/O�ʋL䬣XP�/`|�J�g1�����90�7G;!P N�����#%N7�-�{P&_c�\��p�|β��1�e�Bg_K�k@*@S��k5k�bJT����"+�����-xp�rW0K�q�� �'E���Z����ڑ��S��࿋�3����A
0/�gN6
�s�~�ʇ� �T�+e��yX�=:���&���C{+9)a�&ME��A�p� ��@,�����#a�	~����^"�����0�b]��$5�t�I�q^�����ˑ_�4,�@��q&�{L�����1{yNp�"-���R,�4��^e�ؕ��("�u8pv��0E����ɗ@v�n���y��f?�$W��7x��-��(n6�z�ߴ�ϭ�܄!�[����l�C�ڒ��[^�Y��G<9�:g 3jk�cT��d%��X3�m��M]Pߺ/���d�����9b^���[QU���w��4��	��r�X|B؛�L�]*4A��.�)��W��=U+o#nǸ�?z�)��4�������S�p�ga�z� �ג�%�:Q~o �j���s �,�f�"D�4����p��S�a��dI�l���N���6�~4v��+i���l�ͱ�d;:��jB��0�P��h�6�D�ڌ�ӱ��z7Ě`#�y�j:;��c;���9EU/	-	K��k��91��9u� Q�0�q7@�	E��?&`�ilaD�%��2����[��H�)g�铙��Kǽ[��t)C�ϗ��S�c�d�����ƞ\aw��*����K�s�.����]�a�����	�	����9�u1=-��O �H��2v�_���F#S�	c�[��%T."#�2�v�{:߿��syq�;���9	�[EU���eo���,�����\X�I4��x_�K�Ձ���	�my�Y5B��XY��x�qw6?8�C8�=uF �����j���|_C���_a��D�S�Σ���E�7�r�|��rn�㜻�?a�g�)��E�]��2NAUw[����������3�WӦ���W�檛}�G�mr��7���p��2��mghy5E[	� 5%�!"��}��]�bͫ�.<�}S�5�����-���M:ڿ!�q14�&��
�"�S'UG�.��zwl�n��a�<$d!?#����Y����`z�5����E�����O�j������)���=|S�O{��v��Q������0��u\`�a���/1ȓ�F�y��J����O�rް:E���&�{*�bee���A��窷�B=����6��� ��-����0˥n�-�������Ĩ��KMF?8�C!��S�^�~�Ǒ	L�����둙5�l�l��(��[�M?3Og���[�l��~�wr/F?���D��\M�\,�i�<yZ�=�- �m]�{���p5L嗐:ޔ�ì��88ǘ�ࢧ�*1�%2$��夁S���kl%K:rjqZ�#=�[3`��_VD���ԡ7A|u�����#��Qү�o�]!?YO=��LH���R�7\�3���s��,I��ȕ	N����u���Fo'^��:'����miȎY�?�A�Hݜ
E:���/����q8y��K��.�iW�8C��5�������Wܼ������W��_�x�vǹ���.��ȟ
ʊ�7�F�/s�����\�A�_��V�/�8)c�c�%<��}��@s�S�_����?�aA�T��w��j�X�����9o��>���h3�r|O�Ry󟼳݅��j��x��KF�*�1���n�I,ݿC"�w�jM��KL��1k裠j�%A��| Ճpo���dbbz?a��{��d
'Mu�:�v=-����y�Up���Be���_ǡ��Q�X;gPԐq��9}�t���N1��qȣg@��#�� �E������Zn��=4L�G�z��9z�R;U/"��"=���	��(wFg� ��X�mX|_�6�{��B} #��y���������G�0�cX��p/���Oռ�iܩP�oݥT$����� X�!+�+����qj�4����������1���8�jÚ0�,_"�R���K������^�b�Y'u�6g���d�
+������p��}�Ju�� 'g��+}q����57w�9��(��)!�}/gE��,@�Wa�M��9�(�h����
����mA��PB��.IA:EJ��;	�Nii�.�����f����{ν߿��yD�k���;��c���n�P�V���j|�f�Q�3o��[��n�5Q��)���R��fM.|��=`H��nŘ�t"���4 ��*�|�G��Ls,�>�݋[�7��GQ���*��*�tO�Տ
����|D���K��9/��/�?�`;Ra�'.�P�ޗ�D���iJ�p}������c�_J���-��rw-���sn�T*��z|�[��}9cj����OP�ж繋�Uo�:�8�A��y�İP_)�,"	I]3��4d+�����nA�D�G��X�`tr�����_f��~ڔIs����BY(u�t,�%��Z��m*-�-)�Z~|~ך�H9������U��9�,E>��r8K)>�l��H��Gt�=�L(?!&)�����+P9Ej��,�����tZwF���^��B����A|��P�r��G�����Nd�n}��B�l%֒c߬�;鈙jqFҎ_FOA�E~��cR��x*�~�2b�nt��@�	�N��ӻ���k���X�
zlu�goh�V�A��I����{|e������Ajʾ�D�A�~D3���+M�E�3S����AO���m%�Zƹ����y�U$���ʋ���/7^�"��5 \�!:�*v�C� # �����;�*{V�;��%z�<�i����{�F��0&����E��'KQ"�����r'��1�'^����T���!"�6F����bxg��h�ɿ<Q�9��:�����J��%��X���̋�̋
ĩx���m|i\�G9�+9����ɪ�b�5߬�����OD@_��YJ�1�7��!�W?L�Nի:k	�g"�S�Ey,X7�֝�-�Z�g��;��1)+18��QP�q�^�+��j�\���w��P�O��5�����^��!m;�/,,��N�Y.#]:+'�<�g���I��7eQ�o���������,�0���R��l��`���Y*�F��e���󓮷��Ϲ�;o����p	m�u΍�8�#h�v&8)�����rB��Q��dkR��Sw�D�b������|�jM�Oj:!+�{F�����]��uv�f�_���ʨ��$�`S{d������#�v��X?LF�2�y^�z]�	(����ῂ�-NN$3�S]=}N%V���x� r�h��sN�4p3?h|��P��0恡����!�H�!��K���$�i
�ܝ��]����	�WfL��L�2]�9��=%�R�Z0>)#�R�S��䈼�{П��Bo]%u�Ͱ����8���wS�
��r���(���e$���p'�4oBV�/�X�6̼����{�>���`����6�3��M.���y_Jo�?-TB�1`F}����w�=~�|\q�9�&��B�B�HK�y����w��,>�Ǐ���irˏ{�}��[I���h�ŗ��~P�ex��"�]�����{|}�z]h��55E�o-Z�o�[����C�nP ʫ���Mȣ?iqpz��z��f���hJ�a*r}ٝ��@o���W����r�6m����9
+��)�$c+Ϡٟ�4�5�Va}Bq"��E$��Ե�&jf`�u�;���6ǌ#�SE��v��������l���]J�ٓ���hs^�]ى�Vz��Jd�N:�#�Z�GR�@�Z7�q�}K���������-U�bQz��$>���yK`\=�|w!��?��[/�(������E��S-��H����q���M�.�[Jl��yq�g�m^�xw��rr�l�B)�Q���鞢�ڬY���7?��H}c�U�.�n7ts�%�{з�[���J����b������i~��=�?�ٍ���'�"h�9�����m_�?o�񛴚�tR5�ҼY�i'Y�T��[-a�G�}�{�CN4�y�	��^���0���CAz�l�з[�q�����M�j�0�\䲋�-r1�܁3I�᧔�f�ժg����Ab����x�OH!8~��|�B���Rj]&\>w8ؠ�g��t��L��ֲ�6-����ѦxiQ��o��˺oM��Y#Qb7H�f��y����Ӕ~�k`���&��F�^6���:����#�C� ��- �\T��u��66e�Jq_���|�cT~g_0��}>L�e�*sX�m-4.k%�!����V�f7�l}���	f�ͨqy�����������R�g-�L���d_���˖���|R ��zw#� �y��Qv��]/߅�q�M*'�S����W�d���F�*��_�А.�ݘ��}aƻ6n;}H�����1∯A:@Aam�<́�&�{;tXd�%��s�����{�ƹa���9��X�4�cr�+��e�~�@Zc��ZL�鼝P����}q��;%*5��\:��'�4��*����J�����mٹ�� �t�i=t�_B��*����L����$�����O]q���! !�*$��{�qu�H��&B�sU���|�����V�1���*�l�I܏���_�����zC���S9x��I�����3`�Jy ��V�~ŜL\x���껵�sQF�>���
�P� ��["��i�H@�:@��� ���ok�M�[cߺ	F^(����5��Y�?��D�mlI_�joOw|dܭ��yY��A�[9�nC~�=��R�,��b�rcIf��##8999o4���n�^��o��~��-r3��B�|r;LZ�ݾ�8x[� #��1�#Q���t�*e�_�7��D��Vm9ݽY�'�C�g��+�wǟ�`W��0�o�NTy��s�7jp��`ﭷ��ك�򞅄�9]���b���f�����"[��y�f��ܭ�&{<�J�� ��Z�>�+3�,<!	���ߐL�<=͗?��� b����kk�%�ߩY�(�[���6(��^z��Ͽ<#�G����|�Ԝc�?�������Q���f�?{�6L���ð��
�G�D>��+�Lh�n��ў����֜�s���<�����������0�%>g��V��g�FFjot�`޿�����bB#ꓺ��1y��v1���)?�7x�yx�L�:���������#MM͟�~��L��"�jHd��]P���32Ύbb��>��Dj��֜A$�[j���>|��ya���]�
WW�.���O�s�|��i���QZ���L%�_���\'�*1�7*F�vu�͊:��o���`X�+]#>)�ml���s��X�ak�
��Uצ��T��_g��Fc8-_R����8ߘ3<Os���0�K��_�
6��4���]~+]�hh	oO=���9��G�}�A�n��d5$fܲ�����s��e~���I��-�a�^L��ubb�>�@�/����.$��پ1z����^�����0�!���'��\�x�n�h��x�u��O�ש~m�Zu��gл����&bA/�%�n���ޛn�u������x�� �K#�{W��~��9�� ��)j^��P��^fz�Q� �t`����b�d�$��]�����Ꝁ(��[cI=�>�>�`È���-�\�5�j�u�&�h�߫�y�.�R�������1��0�O~�?�vUa�ɢ�}�l����П|��5$�Y���ǩ���Z����a���l7�Wmyll�1��u���Ʉl&8
/J�B
��K�Z�N
���ОM1�C��8=�N���*�*e@1'66����L~����'����v�d��J��<�9�)�OR�F.�/$��&�2>CF��ZU��;���W�]GE1,��ג�����Vc@qJՍ�i�H��|*�����;ґ�F-6��27���$	�Z_<���r8o�=���L|����)|�O��F���f�ל9��Ny6[^^�ފ%�5)?�իW- ]c��ic�]u�^}�j��9�+�|�	~�E�_A��o�,)�M������'$�N�|9e���C
'�Ϙ:6�V���ԏ3�~Nj�z�Pj>2�'�����5�ϳk��WR�}3��++��J oD�;J���A�+�$�S����
ȗ�ΆJ��û��̓�>Zك[Q�)F�o�ghk{�fl�_�␑��A1��?��)�sl�� nˇD%��Rk��ʒ�͚=���%;�O�.7�D�\Z���A��Cg��q�Z�����̎;��^�_v���~5��n?�����tHuq�s-����2��bTxVkͯ�fه���5���4���ȷ��GR�(�+;�ʕ��(D��1J=��ǲ�g�U�9�.Pl���?$*/�ǆN�~Wk��fY�>��.:����^��F�_Ϭ��Y]�85� W���η�8 \I�,'�Ő#_��j��r��C��-�}����a�=����/F~��Sf�$�~/�y�����; %R��D�qӝ�k�����U��PO�Lb��p�{�wB�J��. v�φ����て�=흃�w���������J?g�н����Sa�a������ѿ,&#V�����0���f, '~}�`�8�)/�8 jV��.>���vz@:���[�{���㷭~�[ʑ
C��'@�P	�?�K?�~Hw}V��k�h�c��zy��u+����c��ϻ��U
TUhq����,��F��oo����$;|�����l����/ip�E��qh�Iݴ|�լP�����z��r����C>
"6iQ���g�q�>G{�w}��u���E����	ԣ1$4t��.ue�;P�!lU�� �F�t�<�u^�FݟU�ޕ~��\��YJϲ�M�_��;} �:d!�k�X�O���:�(
ɓ��A�<(Yf��x�/��Y���ͽ��_���P�����u쫻~\���	��͗GVל�����m-���n���A��������jam9��L�a瘐'���H���5+�{����8&ݎ��@��ϝ��K&��r����[��E��OŰ;�=\��X3���?v�M.��������0�~�հ+4y��Ed�f�'Q]o,-�߾s4 @���
�Yz�1a�� زR�-�XVV���;`�3o )�&�/�Է��㣥:�=ҧ�/O|�O�ؾ��Ea���b>������E��_��ϋ$<A�c���he�F�w�nB��98
�� cvW�%�'�������TH]�|[�\�g�.
:�r�����Df�+��8�<���Ӌ{mn�T�E�{�h��� ������<��x��)诖�ުW�M�� }(��q�?3Z��}|BpWp`����Se��fBwۘ�VU�K		��?��<	��SA�v0�N}���nZ��h���C/����[:�� &o�|�*y�o|���������v��k��_�&���P�w�P�}O�A��@?�,=��V�L��o��m���
-��ܽ��ݰ������`�N�ZX|��s!g{���Н����9%���_�KK�iAؕt%����n���tJ��9I�9%�h%����j� ,�+���f>��ф�����@��L� d��.+$��<3�4A>/�ߺ��m;���QY�FT�ڶn?�Ǘ�$����DD�?s�������KS��/�۽����Ĝ9��Ey���%���>C <,,,��#��O���8��'�ֿ�8��"���� �HuF���>�Ըu�Faq�c�r}�L�n��A�kk9�F�y+����T�ҩ��gAF�m�`C�$��Z�}�{�e{y� �X�`?�DUiSShQ�\����4ϳg�4xxx�/(��� ��o�߷��T���r�IZ7n�6Z�-E��Q_#�[m����]����t�M_όg2d�GV5�s���ǌ��4�+Փ�v_J������������洈�����:�N��d�� ���	߼���,!��ܶ���B��h9�Pp��ÿ�{�N�5�j�-�?m��\ku ��Ѩѳ�S��v6���fG��l?��M�ɻ��ܚ�U������ 
�dg��1���U�������-7���U�Tj�M�u�[���brb2�'l}��4���X�z0�����8�U�i*
�~n5e�L��NQQ
7��z��@�؂ss��7
뛛�e֩��J�'-�)��󥷶����o	�>ʮ
TN�9ٕ�v`�sKQI��n�<k���՗���oa�3��	yƅ��Yx��Pi�t����S�j�;m�#�Ù�����.�_���hj$�ߓ�����}��2>!Q4+���s)�#-����P}��OB����߀m���F�to�ȕ��)i<J�㩬�;���C�������/��mm����]����������qX��dd%K����?�����PTW'w�D��4?�V`��CS3��Ǆ����~U�|/<�c��������O�C����WQS3�np��G�k�4��"Џ�m�"3��~��
oߔl%���9(���f
N�:X�'�:ɼ�m�)#^�4y���G�%`�:9�AEE]��^�O�%l��IIIQ��4{ Z�{=��?<x'[DE���ӿ��$#*ټ�֯N����0P�]���c�����[Ӎ�/� {�ʃ��\t�grnd�r�p�y�U]�o�-0g��2F��R�ƠWg�ƿ�"<�~�ܜ�Jf2a�	U(�
ϡ�)�����PM�u�]xś2���DEQ�I��|��pܤ,���F]�x�]S��t`i�OI�x�����)�ŭi�&czP�����"y,wE����q2�є���#yʶ�Z��5��tt��ө��V9Q�׸O9��jsE��%�ћ����>o~?Ӆ�6������7_�iV�+��޾�N�R���.7p��Y9��~���� 	���ò�e����'�t��̀n�B@�~j!�4�V���@ �?%��Tڰ��%TǪ��c��PV��roB"��%�~�k�vQ�3���&�(���r�9�f�Ak��/G�N$��y={��|�w�;"�38������d�C�{ֲt��d�"�^2u-��55�D��n��L�K�s�ԁ[�����(=���[���hQ��F��ߤ� !qty�sN�+ǯ���|�<�R��ow��m-ҾB�A>�^�,۶�P�Ϯ��p�l���)tT����~���P�Mm���D!/O;v..��4�XFĚ�ģ��=����8Y8>UD���}��k.�+h^���e�9�Ɉ��]+�<i��:�%P�X3��F�"g�P������r*��6�2GX����fҤ%p<�����U�Mî����{���Q�ǋ�C�_I^���*�����!�V�i��h���kn����ds�d����,X�h���_���I��z�óU�`�\��X�9�mS� �����T;*�A����*2ى7J���ZT����@ l����/ϏW���ע%�N�`]�E��hh��Pě�������-Gd���^?�j��~v
>�6yN���Z�KRN�i7h�T����]tvvF/)Stx�W^�u�v��4���o���
u���F؟e;��{����B� WLMMm9w�.���J�̛�U44X,�?uHj�����o� �W�V��`vS�oh��Xt*Z����^�xdU���a�1;��ym�+Jy��T$ZK)��P�9`��[p�J=M�$�Ϻ�}>Ł����Y{����3=%��Ca�@y�������Z��,���MoOՏNM�T�j3�-��$!~�ў�j��hOF�d�c�<Y:��8h��p��6���m�&��B4��G�{��6t5��1:&��5���gN��w�c���k	d~u@��p��Ҷ~
Ec�]���.�99QQQ����f��!�U�/_f��d2�"[o�x p%����@��F�s*�L�#�'����4!�p�C�yu��m��e��$��n����wX�I��ן��vAi��,MEZ�C>b�Ps$38�(޳s���1̎����
��:�I��x>�b�Jy#�yϵG�h���b�P.H�u.���p�����T�[�⺍�j��Gͩ�KG���N��^��Ed�	���k�����Fv�%�Y���Ծ9 �LMT��o�6@ܤ�ك.��W,��0+v���Q~N���1��/�&F{]�o����p��&����G��s�	�'���:6�ݎ�<���ۡ��#�
PJ��$4:���A�p���z~Pf�)��c���f#��&��/��>)�`�=�|���)��r����u{��PY�j6V���1N�Bg����|��]���ڭ
�������I�z��ı�8�ס����D���ͼ˞�z��������^FO�I��pbB
Vt=��&���H�_ϋ���􈃟���̵`A�HSSS.	k����<���9I���==�	C�R�{���DYR�~��3����-���xH���Ϗ��@Hٝ��V��(-�N�O1�<�$.��&�sMM>3K���z��X����.f�+�b��N��<6�o�ҝ�Bw^@7�A�i�e�U�L�������{���+tbד�����S��4uX��C�A�\n�AUTW2̢||dr2�Œ���FL�N����w�J�c�<�",�����Q��o	��C~f��g�xA+�Z�3I�lb�Ka̰:5�1���8qC%X��絍���cR�ۄd�?)v�n,��,^��,i9���o"Oe4K�Y�a�QTEE0��6 ""RQV#�����Dz�g��$�|UUUt?�Opʀʟ�ϾQ��%�P�^z'm�i��^�zt���G��i׿�7_Psf-.~�l}��4��2�G�g{�Kc���h���/�k+� ~;FE��S��ϡ鵍�њ])�nk�Z�3�?�a/��� ?��r��A�+ �!�556��+'g��T��-~���s:)++�����%�;���1�]�#�u�zrkd���Z���_&����Y"zAɓ��0q�m��E�v���P9z���t����z~�3��Sn�v�E��`��t?�R�S�9�\�PK&�%%��I������$���=��嘘<J�Q(�z�$�<k��rHN�h����
�������*��i�-�%�c7�^^ƀ�ë��� U���hm/peI=��
''�Tn���9y'�,�a&�0�AU=�b�����zw���|���\�t��7�Z���"Ǹ�^d��u>���?���p��9󃠤�ht}���ŭ� 2P�T�B�aP1:�S"@۠n���5/릅rD#^Sa�����J��ċ����tGC����ń%�Zg7!���m������2M�F�"S�z��:5��7��ǽm�NiF#����m&e�F-o-��qu}�Wx���M_vrHH�1�y bҭٞB=�����b��.ڌ�cړt3_+�}N�hEhY�h�$�W*��g��:|��k���^j�8��c���0�/��'p��M��C3�!S�+��J�#�(�zkG1�Q�xB��Hm�E�khIO�c�-�R���լf���m�\����>��s=]��'����`��U;U����ή?�~i���(L7���|1 ;�^/��E�g�p�O��8o꨺�X(Y����*�� P�?�z���E�V�҂��L����>u��։(����%%+#c���!����os��KaG$
;����u�M�����ɒ�@*S��c�˘�i��^��mtW���8�~Kq=*)�$r�$q���F�,�<Qm��O�D����O� ��0Κ{P7e9:2b�~��S�h/�¾a<�4�(��U�fRƙ|OA�cS7r��+Xu��R>��B1�4~h(㏊�yyRrF���0~RX��c�L�(<D����ol��6�½۱��&U����G�����:�	i�P�n`�����W��Z�0w�ɕ�R0������ԋ��vӁI�)Uf$��x����L�d��h�=��	��ѥ��K�����k|B�n���Im���+�H�9ئ1p�o~P�rG����F����B#�\0Kv@��f|(��Uǵ�H:!��{��2���ɪ�|�SA����}�2r��-��i�B�_
e��T<%t.R#�_��%Y�I��u��PZ�%�� ����=��t�?�n�j��s!��J��Ǭa�j0|@����<�=�3ك���r���ɩ��a���<P��q��-+�[;����h����
��t�����j���^"�PR�d���diZ���O^��L�z�^NXޞ�5>>Um��M�b&�U/�gB�v�׈������u�p��X����<�X�4IrW�bb���J����T75	f��x����53�B��h�c+�N{���cC���-��ص�\&_�9²Z3N�1��~��A�N�ӧO./4��9���cc9��v3߅�J�o�N7���re�|�t�u7�um����8��:z��[K�<wI���e���K��rD��fv�Y�03�:�b��SP���'���u�iG��= �G�~A���8Ƿj�CuTU��'���m�N&ܟX��Z9v�с$):3��d�s�6��$I#?�?��]�>���ߨL�Wײ�S+|�n�۵D;3<e	�8=���GDBͫ�nE*�c"w~f���lT���}]��D��4G���+�uf�6��:�������.d�����j[���;������c>���,.fAe$Ń�����6ϔ(�ʥx<�?vs������,	 6 �R�g��B�?�J��m;J�j����ōG��FUm��]dx�8��W������f
�V��P�w��u�b�qGP�7�=<�+T��H��ίG�'FB�b�ފ�ۚ�M��f(!Ǳ�?��쥤��U[�^h(V_�G�G% �?9y~II5o�>�J&W�<[�ccc���ܙIN���nz}��n������/៊���(��,%.�%�P�}�P[{�f�A��_����RRW�մ������4�x����p��~}���Ծ�Nz�[��e���=$or�Z��N&'[�Xh6�L�!��D.sd 
.�&��*�)ccE�����F��~4�e,}�x�\�20�t��B�f�<'���G�>{�5�ړ=h(N8B�ɸ��'᨞��V'�!�[�����R�Jt���/�r2�+�����&�<�)��D��|0]4 gjT�ֶ$�����Y�0_]�3��$��$�?��Т���- ��@}�F�u-�-vF��ʚ�n*݋o6��U�O��p��%Ѫ�Z92�{��'��-�^?�Ǎ0}64Ð��˜���2\�;�?p���"�-�&&&,���J�װ�]p���J���>���A�Z���S1��R��Me�館4������ 5�#ZK�߳�{��� O����t3Z���`����ju�8�����q`�;�.+�Nr9`�����r�0"]��!��y:mҒ���BA}�q(�̿h�D���~�}=��Uo������E�Lj�K0�2�{0'�1
�G6�e�a�b��n%�^W.��=HLNN޿��w���y.��\��-%ؙ���:c2T�4�~���`����u���(-gy��Hz8��r}��(^$��c�d�l|����oky�VW8/�o���~JA��^�\> Y�
֒��v�ڑC{_�5�rٿJެ�e���&�u�V9n�����v�ceu5�c�%e�����ˣ	�y��A/P��Ō�#?��hN��G�;sGm���� !�}S����������saBN��<d�Q���{�o�A`j�~��h���B@@`}s�w<R�(NR��w�����xy�9�M��#hj2W�����{�{���?��) ��~����a?-ud5x�o��3Ivǹ���K��5fe�0��)Ǥ�B��A�	l�Cm]��f��oB����S�Ǹ������g+P9uo����ļmq�=5���޲㌣?J�>�%%�P��d�3`m�&�S��5{�����V��"A�vU*jk?���J"NEB�~12hu`DTY=���F��CRN��eC�&�$Y�S���mm�����=X8��<�0�3W���X�
>_�ݳ�s[,�w
��@0������ث�e��v}(r> ӳݎ�� ����F��2�r����P�����&SC�}y3jy4�h�~f�'>ઈ��ENC~�TF�2�r�]�����ӽt
�C��p2n�Z����@�ä��$���UϷ]#�{6��Z-�p��+��KX6�	�	�p୭H-�_Y�f�:��a�J�d������?磀'���D�����T	#�������8-�J�:m��:N׶���܁����W�U�i�e��E���:M����?���*���!��V�I=���VvSSh+�Ϯ��	0�H�S���{���9���SQ]�e)z�0��5���lg�ˉ���	2��6Mu怭6�E2��4��c�BJ^�~�a��f�Roj�aKޠ��*��/���M������,��x!����9�{~�� ���p\�WݬJ�Z�x�f����É�LQ��kd�3�71�����K�l�N��P�BhGF��X�\ҋ�~'б��2��EB��_r|E�Y�W��#�0�����^Aq]~��5�d�hǧGT)��m��������s&1lx���<�d6ڐi��h�t[��C6 ����	k�|4,c����+	7'��x47j-�y
n���8�"t�%��0���
,���Z�L�X��vz��u(���\���q���g{ˀQ�*=����������^2��5������sv�k�ܶ�]��ܯ����зڷ�;���&����!���ʑ����Gl����ʰ�k�\B�%��y��+�jj�P�R�rM�l{8ƣ��5��~����]��|���v~�n9�k`T�����`�}���*�O%q�(�.�z���ߟ�O�1�e�u?�
�ݩ���� \��b����`3�l^圈؈�%�W�t�_?�d�>�w��������h��s�-�ɼ����	�P���s�ig
�=��ˤ�(��S�'���l�Ar��7r^�l7����ѽEù�	Y�;ѿ��BP��HND?�n�y�ɮa���X,����Ƴ�	b�VvY��ᢹ`\U���o��'�k*'_�ɗ���H4�9y�wY��r���K�u��Db�zX������ݻ�h����&������[��:Y�e�D`_�b��M�K�0����_ǋ��L�
HH�w����"��:osLY��/쏞$#܈HJ��3�<�z(T�5DL��Ie[x�v�&�x2�8���s��J���yyP��z � S-}�I��EI�U�e���{[�:+�׆��V��W���&��,Yw*W�ṠJÓG?�h#�ĕ��A�r�&\�d�dڪ������ o6K��~6���K+�$�P�[��W���<1����X �K�o�w��*���*v�����8�S�(ZJ��Cq8��o��~!}��H����-�Fhn��֣1E��G̓OdP.[��Ժ������������}N����ꂪ*��q�Յ 	%��rF%�`]t��蔡�ў��J �?+EQH�%w�L�q�'�)�9�%M�Q��d]B�8�:�9l�uY�:���o9iV�a�3�T7!>��&G���g�j���(�9`k�?@��%)o_���=�NV��s�o�|K }�,�`C����lc���x@�C�h<׿�˅M"�l�z�2ɹ������)K�u�76~�҈�kT`A[��&��[[}�ǡ��>^O��'(�eߣC�eX1��w�7ӣ?%IRyw�?��%��sQ7�Q$�ht�Ӵ<>����#�����]��p�n>�����"��vގ�n�ԍ?<-�����̫���":D��F�4�����J@T�$�)����"i���%�L���$O/���ᛤ	ֲ���._��n����Q�%ȷ�����]�~��b����_��ղ�e-I��t��,��~�9�W,u.�{�9'�\O��>̷I��?��ke��}u���_j<H�qT�6
��>�C����^'萴K�a��0O�Ϋmń<�9�H
�4�zU�ʶ�J�����H�y41������)/���6���o�N]/��h�8�B��9^}m�a_2x�F��N�
)w�pdQQQ���������
�\Ff2~>n&v�I��a�C�=[u�7�3��Qo/�	��]��?|�-�cX>n�U�1�c wL�TXc^c����X5V [?��	����\�,VɌO4ҫ��h:���3��C��
&�F_6�����O��0(�g���H�ݮo����ڴNz�<֯WbCJsr�}���/�����@���+{��n�.�:(�	�M�~#QQ�9����ϧ�$��V����x�g�E�^[��M�<)r�?(�wZ0{�s`�G�PcyW��	`����.n+2��C���$i�w�r�D��7���3���#6v�<,%�z%bz�ֹz>�ny	�%OM�1ߵ���J��X�᷑��y�d���i7J�J"�8r�(A�e%z�� �t�t��c��dq!&�BͅQ3��������Q���YIcU��|�H����e�Rc�ӗ�'n;*�/�G��Γa��k��-�:VV�/]����)�$���������j�c(�j{�z�g[?�_XX�������I�ˍ����,\^6�I��{]�U����h�d�3�%A���U+����c.���k�%�����^#�̗L��]
X:%P/�u�G�?\�ݵn{]K���s�c��{̲φ�E���.�����;X(�Z:D�=��3��I�L�r��]ԥ��Pߛh��ҔV.y��q�:���ڭt[
i?�
�W~v�; n��)ϫj�%�ĉ���I���$/�5�'������n����m�F{��POBuu�Yk|� Ql������W��Q���i����t�c�H�F�J��;��$K�!�"�EJ��妛[ x�ё#X�Xg�b����Ԕ��qx_��V�"������K�SҰ���F$=j�qY�NfQ����� ��8-��;��[0�-�l��,�R��̲L�@��>j�R���c?*mQ���#p�߯AϞ0��H\Y�k���_4=0�@t
�z�M�px��^y:Qux'�La���{�8Tj#�\D9B�耹�98�l��q([	�~������c
��FEk�~�Bc�^9���>��i�,� u�}�����A��ô�Z�q�{
9@�fB�+�b�-{��n��`2�?�K��S^����H�9�	��`�]@$�p��p�T��t[�$�Q2[�٩�`�B��
m�#�t}�<��/��o�5�X����a�s)?�i�
����g���2{�i��zT?���08����d��y-�ԋG���@.���u��,sG�a�G�������V���:~�1������X����e`��<��	���@3��R�յr �y/��y�XHb"QeE��� �0�rG�$�ϭv���Y�|`������TfNw�r'����,��G��Ρ���MW2Rr�����G�u��l_����j1���e�Z��T]����t>z^T�0Tqh^T[�3))	#Y�H:w�W�A���Lɯ_���E�������#^�X������ⲥ��Cs��7�`����$�/q���غ+���Y�qε�J�,ĺ��q0;N��y���`�� �}��S/�`�K��U)��+�i�׭��l�9��5EO�d����W�<�{�zu��n'���A�Ļ��]�I>���>�ʵ��"w���B��b�o	ah)�YAhKM�H�PV��u"����"2rl�vC��X�w	��/���qh(��ȓO!!8���sAt�za9V�I�!�i��6����Nua=۩gy�~������'�ڞ1�,��X���1$���!��uo6Ԛ�b֭E��y��҆Vل�at(���朣Sj�;ZFE�{M��.%�H�<i��{�S��<R�ؔM��]q��\�E�\ta�_B�/�\�-O:�F�-\^��kYzU�[lI� �7|-�iZ����RdT�4j����	ͯzyU��J^)� L#+SSZ�����\I�Ѡ�^���ia�/9'+k��?*��xsr�9_��H.��x6/� C�g	9߇�Hc�8i�� F&3�}\˳��2���t��ȋX���l�d�I��e��ȝ�-����PH>;�nf8`�M��M�eΜ|���?��`8^۴�Q�Ӕ�CH� ���p��I�����v�����E���eSy��us'�	lfp�ɣ����y2G��J���_�����6�FF�
v��Sሂb� ���am�4�V�Ы��C#��^,��D2�]�A�<,��&��x:Τ_^�a�k��]�4����\�2���ܴ�Y��?��o8:��04�������*?|^�Ѻ��:e�,�,���r ���T_@D!��,@�G%����]6AB�3`c�ZO-�#08��,:�#������c�T�.����Z<���s��kC����֥PCi U��-�^�;�B��b�����e�ٸ�'�Q����]��6[��Q��,ź����6d�W�3F�T]���]���ְ��̏��6*N�fT��5H�
~�Y�[��W�L�\��
"&�b&`�v���^^�o4���(��߿�u��907�����W�(������
�ngg��6�c߿pL+�NN��-;�6K�J.b�eK�>'��G߮���o�u��[��^���6�=+�������<�^|)���j?�N��9D��a��-��������zi�1xy�d�Gɱ��Q��lV��ٖ����ؚ�~y�z�P�9����Pd���Cd�k��W��l��T�K�8�x�m�&�9�p���A;��*^��,��ҲX�$���>Ȅz8�0�ٖ2-e��RA�A��]+c�5ȥ����$y�L�iK���(X3��L�(>�`�h����~���)y��EEE�Ke�*i���+"22��v2�ttV�2�q<Uw�k�U��X9�{W��C���5�$���Jt��s�c��梯;4�c�.�����仜w��J��~[o�2�Rf�~|i���u�{�4�-���U��q�w�{֟��h��(4B�T��0TA��^)�k0�};��]��3���y��C,��m�삂�t%J\��m|���Rmm�֏�]�fݪ4��پ�(T���5���YR���ln7/_�s��y:
��*&X�\��j&�HF!��+�؜�r��`(���ϩ:\��ٝS��C%�y.+.�U�m����.��Q��A�/C�c���D���ySc7�s{�KW���!����ŏ!�ێ��N]{O��t p��zF�B�H>��3�׾a���m���;a'f�yď��X���1G�r�ix(Ǒb�$�����Fm'�S�U�\���&��WWÇ�z]'�~��Bk��|�)���p8���c�A��;��y����������ߟ���:7ȱ=x��wc��;J�0��q6/��QX�f�.���U�L�y^�7+$e;2��G�[@Eټq�4H� ���tw(H7H�K�tHwK�"�t�"�"���]�����Ι{8gٝ�����uϘɶ�E���\{�}�7�4Y���o�o�;�9��]���Gy� �B��ɭ�i�� p:	�G��Ղ��L	]�csu����MM�"�����\��^�Wb0���Ƨ)�Z�P��|g��x��o�F�9�,V�ڑ�����{��ԯ|��S<��orF{����A�+��^���SMM��S:B��)��px�M�*X���Z�TdR�����I8�kR�rL$�'j:��U+K��e�d|�}{��2,i��÷o�*�5�x򦿫6y���:\��uQ%��=��OÆ�5��]O]�����T++�U������]������UW��zZ��B ��ϗ����"c����Zb��ML�0��⣣�_��LxR�O���в�7e)�����r;$�Ǌ&�����i�2=+>֞:9;������#Z���  \�d��'�n�����u+�����N����G)����������z�����P�u{�<e�9�Q���NMܼn�R��m+M��M��a���"n�z��x��Fa��F,ӂ�����D��M���#�Oƪ�E>�F9����4�j��Q&�u�Tk&�ͫئ����T�N���Vk=Ѱ_RR�jP³L<L�ə�"={�E �K�{�"0a�=���n�5`�LMԎ}����2=�~��@F���x ��\ӵ׵�w��ATE��� �%�Fֈ{�B)�?W*;���K�V���/�6��M����SN.ZԿ(t֦�L��]�E8s�[�iH����]b{�kH2:
�m$��I�foZUJ�h�Ij���G3����K��M5�Q��yٲ� �Ju��e4[���",#J�x���vc1{@�6�ʜܲ� �;���-��{f�-R¥�[/�L�]d����|���[�:����02�Ҥ߼W�r~��[����U f�
1z����F_�֫!�=J�-=!G��u����Ϻ&�	ϯ���TÉ��'��!OW[���}p�A� ��	䲠�M����c\B��ť�����a��z�7�3�[qC�/�D��R(�x�:�$s����tx�Ջ}�(d�B��d���q���8���ʭe�������u�v]]lS�m&7<���W@I5ߟ��W�'��Σz(z<eR-�|����)��\�<��������������ޮ(o���[�)u���cqy{�����=t���l��9$0����5��WR��3G~S���Ho�{�LpK�b��Ȩ:z�~9cE����*���ɿU��Ըc�Z����7SJs�_�GӢ6��n,�O��!�N#�ɘ�.�!�e��?[4$���9;]����M!x��~��X�Os��`�5F>�Kz��'�e�^Ђ�Tc����x���Oy���mf�S�2��ܟԒ�����3�4@�Gɱ[�$f���ϒ��ۂ
��"��[-\	���\�~Ϯx�R][����o_�� +r���1��_���*;��la����{Gr#[�Q"�����vѥ��h6�����#|w���"'ǲW��,������ �Xd�V&&�kڟ>�e*�V��������K��J��XM�yg�ۨ|������B�Q����Յ����~WW�f�x��/R�gL�lYF�X���'�'E�p=�*�W>c���fs�{�&#?��$Q��N�Z~嫝���N����k�֐︕z����T�8LhV˲a��]�_
k%�vB�Uz��
:���,p+7J|sx��t�� �ַ�1/�sǽP���sU��������[��O�j��_I���]a��=Le}�gN�?L�T+RCdrg�y�������_��Ԓ�H����VT(�
�E�ک���lq� 	1���ַ���w]t�V�!E���p���8d�~���������Q�:�<�l�����enn���"U���z�!:&f��[Hy9��V�X���d��(((t@��c�~�����p7��a%��Z�MS8ꦭ���z��H���:4�imS���W�o@��0�}�qwuq�N��O��	*���i�
X��+a�	�1C�.f�3�,����?��ba��L�]��T�z^�Z�����"*� p�{j*��@��T�5><�Z�0��q�( �
��^�}�����w��4��-n[������xDRo�\���|��*S��L� �9<��e�X��s֢Y#G2�]"�R����f�k�z��ב6�Z�Q^P��I����װg<c(E<��f� ���]�����f�8�k{�B5��>�j_��vfQ�@u �,L�a�'Kv/R���p���q�HYۮ���ͥ0����7�ګ���LݎV|�{�;T*99�x
���i>�!s��H%�~(��iJ�/<k�V�e����MX��.r9���G����֮D�_��͵��+m���A��&��k7�M�벏�B�� �ʣȷ��DO�{�U��	n�׎�ɝ�l�ií5��,~|Vũp���ם$�����������[WL���_k���L͵[��O[l5�2�Gs܊�����S*@\v��ŴQ�D��Q9��,]ڈ�F�����xȥ���K�l�Ҩ�����G8�1:?~`o�w2<�?�{��W���N�ͶKۑ��N�Q�1��7�3't��^S0�Y�
��[��-��ބ����"��f����i�QJa>�h��P���I����v1gљťҵ�G��1�����?<E���$x��}N�-dn��'Уۻ煌�m�~��?����΀��u�~�������l�h���K,��`X}.&!E}Gd|�Z22���O�>w��#�Sg�Oj��l�Tppu\/��^���\�q|�z�^�$j��sI�O8��ށ�Nv�tb�<�O+�u�6�+�.���>���?�lM�\vJT0���Kl��mg<%yS�TaV���w���@���ˁ�ҵpip�; �?owkhY�bf��kh���N�Rl`)Y�i*����eo~^���GŌ� ��E^,�UU-�Ga�ށH��%��t�b#���U�����{#Y+I>�֤]ta%�T���9�tr#���3e�D���Z~C`3X^ET����a��F�:���� ���zd7<����6���ԛa*m��k�|�Uz�Ӽӂ�|!�A������YvwZ$�uw��L�C��yC�ի���k2���=��i��m�͙t��3��;K7#�N:[,MC\�؇\�d�j��/Hd�>.T��^���f��Ȩb``���������0`�c���@`=�>^V��y>�-�\0�-�)ɲ�I0��9��$-$��ejxz�_�����w;�c1aG:l�zT�?�����-?����S�S�xΩ�Kn�(����y}�¼�:��{�gHhf���:&�
|J�釣,�FN���CL�ﶆƇ��*R��nw�۪���r��]�BԊ1�2���A��?�*uO_��L�_�2���a��lU�ҟݒ;���k��u~�ʪ��a��ɗO�Ƌ��(Q("��_��n�H�P���lL0���,rA@�8�2�P�7ӰcN�RM&
k���.w��Jc5b �Յi0�K��v�e��0y��"z�ud�8͇��>�]e8��T���=�;obf�$�R7x����c;EMd�C�q�T�v�Hz�,��X���p�ZׂR�����)C�n����բ�֬3�j���Y�w��^���T�l���'w�t�����ǵ쯇j(e~{��im��+���@h��/3T�IIH��z�"N��U�9'�KS7Q�Z8�<�^�
�յٳG�|Zy�f�4��z���!�s�`�w=b;E�-���?�8J���������kz�д��[��A������piH}�t�3~������	��5>O�^u:O��]�Fx���U��$b�,3YJ�,�_��[:�ߣ��ݮ���R�k�A
�ܭ�eCp^8	}N�������MMX�Iz?a<	mK����+�-�t�r�%I$P��2q��ڡ^af��$1��L9$�K�N�5 �9U�VeU�m��O<�����o��a�
P9ac��{�~`"U�R署��0!h~qR"��#�~����V�.S�\�r����b����O��%1�@�oUUx���"W��U �,��=GG	j��yk�qMމQ��9E��k$3--�?��{	�E�h���i��$G���� =Y�)sp�}�H�����x�]���K9���q$�߽�����GO��M��JkR~b�}���i���t� �V��̘%���?��6$>�D��6�������j�� r؟y�� 2�#�*"P�9���G��v+��B��؇Ł OU��(����N���c�Z��*����P,�="_>>�f�;�8^K�?���]&2���0���NQZDo�z�N}4z|���;��$�j]�S��~Z�MO~o�j��q=�Š%e�.v�X���0��~������,#�.i�/�*]rK�Y�Zy�G��}=��cf�7�o���А��4*<�c�1^�d� ��wq�k�����+ה�qg�Z^�YQZc
p�'�d�
�hQ����ػ mˆ@fj,qΙ�7/<i��-E9G�:�c�?�)��÷�a:ޘN�١�\��g���=h��f�قV
�>ڃx�h;|n�S+XlA�M�qT�M�����ݑ��W���i��18p�Ә���͘j�[z���e�?�|�cy��j��Q�uj����WF����ă�@�,0���&���S1-�Ϻ��{���a�O�����!�h9ҿ�Z)��ـ'*�����4dv���k���h	��x�e�Ǚv�n��n=2&������A��f-���~[�\���d����?�[�߄�#fe�R�������-h;Ƚ�o��/A���"��~p'L �fL��&�H���@����gv�*����CP��/ם��>/8tam�7gZs��	猦ډg2}�R�@����/����p��(1lj���}�Դ�F�Wh�M�P?�Xy296j�!;6�h�A����U�n�Ջc�FG����|�wf����5Ͷ�ca��n�>.҄^������7�6���Է��Än���j��]�FM�6�X�:Ժ�s�A�Q#zBBC��
�`Q��D�jX��[8�kM*++� ������P ���W�lZNEOxB���(�Q	��;�t7�sR�2k.�Ӯ폂܊\�35�A�[]i\���5�~ch�J�h��̠��D;GqѨ��A�N�Nw�c�zSPh��d]�t��O�Oǹ+VX�m�>�����a�铻/
��؄�?��B�H�3^5s���q+,zW�a.cڤ�]�>�Ƙ�n�鹈�H��tQ�O�7Ci\�|�.�IIIK�zqey鳙V���ҸHh&��V��@"���愤�������N<��5���ɒ�'�o��f�@CB &&���I� _�;�Ķ�嬤�X�2vG�/���E���3y��.[ޗ��/�ڒ���,:�S����`>\�,e�~��aa�l�X�~%��Ĳ�H���ܮ�=��vz�N�VVV������K�g�ܼ��>D N-δ/]�)�zcK�z|5�$�G-jdL�����H�e_���E��#|h:<��O�:��Z&����j[��[��8^����E����,�Ê��[Ea8lW����k1�X��h�󛶥�M^�[���#��:�g�Z/����7���޴�Tk>-��������T�>�r���}�%�_�\�Ч��r�LI�_=>>ZS��������c���28�g�Ib�Ј�Z����\�����,�����v6o��L��bF�d�Fv����j̜�k"O���z��q���Y��@"#o<����C��yy��{{M���KQ��^���{	3��m^�f6�$�u�*O�ﾚ�(���o�g�T��M@�s� �E�������8g`�݊_tz��R7���J��OJ�+���a�9�������U�&��ƭo�h"�Hj\�94���"�هP�X�#��^TTG���:;]Q\�������$��J-i�W���݋P*��{p =`�T���gu�������~t��:�7��Gz<�NB���cY�.����w�rvWlEֶ��Tf�lw���J����~+-!e�sVl\�FĔ��M��z�Lm%]����^�YLU�%�e�e)@!!�.�lV���9�]`��+���y�y�j��_��=j�뽠���e���xx�E��|�y��x�������j�K�����$�,���"���O�v(k2���ۈӈt����<|�r�� ƺ��B�2��G~,��|�v4���$�0oߎ%��)�!{��_%@G�w��(p)�5�H>�����O�~��U�����:ɿ����؃�8�bw��R��]�=Q@�N�?��S�J{_�%,�{�yOƫ$ؐkK"\R.y��R�x�6O��>�.t�H%�5d�ϡQ=�ss��%�><iu�}����YJ�����`��r�y��O�tJ$�v�r��8�,���6�WȠ��w[�6�7��6������#:�`q]`�ND3��e SWͶM/�W�h"x�U��$ �n0]�����������+g7��/J���j�"��>0��pĽx��ɋ�`���0K\\ ��Hj�����'4����|�g��ʚ~rlaJrQob�		)eOA[��xvd͐^������6�6�O^k_$Z���-jv�ʹ%�4lĴ`�5�{���?��tMeEK�PD>=f����c�<��2` ��8c�r��'�.'���#g)�����Y����F)ܱ�&t^��]��0څ�)	��b34}����.����gb����`�P�/��D�����7n����P�@I����Ns���e�؇u��W��\cI�~3d/�����Z-D���@�¼X��T�#��#YB��?�Kh��.p����nE�f�M�"R~�-��P�Yt�)*�[G��:�R~�	-���[#A~u����̜�6�:�����T~�$);w��p춠��X�˪�I�TK�9������g�qW)�{�K^�%QϮzc�)����w�Oʘ�$	���	�q��桡ܸ��^DˎON+f�v��޿K0��*V?	��ڞ�.:�2����:Rs�:,�,����B�3P�]iiSS��n�ᦽ1�J%��u�z:��N��퍕��R�?L�=�_D�+��a��~�zS����KR1{:���[ڴJ�y�9���BD�pp��%^ԑ���Ͷ�����!7��l�x�t7A������?��ц_��L���(���%��-����������lU;:����7�BJM����hU��޵cOh# \ �|Ê��w��'��Q��Nҁ�KYB�i��a�^���fl_�����^BCC*VG���� ?��E��T����B9�M��]��~J�������{�n�bu��f#����Z��o��|�t��$x��왽=�m9>U'�Ѿ^�j��4-�U�����^����nl��<�U��rd���.�}V�Wy���&9k���K�+K����Q��&�'�����gK�?n�q����@$x�a�g��?h�������qI7+B�J*�Gk��>�E��<Z���F���.B7�$�9p[�X�v�	?��^�Q�򥣴n��G\��Y��;T�6Cć	�kS�Vچt�A���L�K���G� �kC=y�Ҕ�&�#^��KI!��9o<髠�Ɍ}4�]��7n62�Y��~��2S���n�y./|� �1`ط"&܍b~�7�i��D���c���%�����e�غ8?/�9����<S�t�R�j!e��'�#�
ITS�L݉��Z^�I�S�'�7��Ȼ��"I��5�
�ف��E'j���u��c�	c�t�����&�ol�� �@N#c��LB\3T��|����D�����A�(�7l�x1�յ�2�f��Nh���ZP�^�5�U-�ʞ����y�k�*;B���NGS�
�Ю1W��h}6�i�i�ơ��6t@X�>�Up`e;Uک��	�F�N�[1l�O��O�l�{b��;�tB荈�gr���}?��Ղ�K��):k��4��E����O��b�",�s�)<Ї��^!d���=�Y�P�c�v�)E�.�q�Q�>�]�������jJ?0�3�+I�Z˽�I-Y���ngx�@���g�"��dW�Q��5(n���A�o�d��(C��_/�Og�dg"#�Ƅ4��<�i<�ͥ��j�Z��	�Hq[�ϊƻ�]!D&���d'9�����e{�مմS<�e���<i���ߠs������D߼��_8�>w�49�����gU�-�L+���F����<I�Tǧ��@�y������Y�A��,�~�^����M�vf~n����z��-�w|C�˽M
yG�ߍW�`���8��C��gf~kߝ�ZeA@����
+PV!��O�q�_��ު>�u��X���g:�����y]ϚB��D���-.t;g"�-���!bf��m:N�B�j�mצ���L���Y���5]�n�'�8ł
�g��f�gp>>>ڵV���ŏ?�kL��y ��G<���cD��Di�s��*�Ol�ZԯO�,)Ը6Q�U{W*	���)��`��*;�s0��W.<���aV-((p��ۻ��7_#[/q9�Y3�YH�SaJc����Y�怨X:��)i�
�Ɔ��>�pL��ts=��sJ��gCv���j"��({ݻ�~h��{�}iHqsy�>������nV��~��+��{T�a_̆�x�JӮf�_���,�}!�)�R�h�7H��V�6�7#�<PX�kC.d���[JV"i�*�~�☥-d�R�oޠ�X���(�u�,[� Mb�JH�ݽarcH^Q�G�7y�S��;�Ʉ���g>�$��r�)�+�|"�1�3e����(?��Y�{�??�I��[��F�r4�; u`���A�0p�F�&�fJ�l�6 �g���u��~�mO{�Qa�S��D�~���]t�cZ��c���I<�w�@�nP�����+NrZc>�nP����r�=�x��I�=��j=�u�xSY�;���>�X<*� &B�p�y��.�Vр��7I��&����8��(Q}� ���v����t ��:��h��N� ���(��I�bfA#��j�'7�P���N��D�[ ���� C�y�q�Ix�Ȑ�xJnR>! �śڳ�ꌿL/�I{o�p{�в���e���0�v���Ne���1$��*��)�^w�N_�Rs7�E��>��o85:���~?T�ڿ�S"���ykDFK+u�\噖���J�O	������5��u|D��W����@W�|����~S+�V�_M��?�i���R]�;z�\�^��N�^�q�K"��r�tΧ����	��lX�їH�]�{���L��@�7��w���nݳL+��l|>�*d><,*�}ቶ`ta�����[C��I<�w	���5Xc<���<�_�%F-sm�-P����% �8��p�;yR��`�j>��Ɯ6O��8�j<�f	q�A���ay!��E�9�e����PM-1w+?I��������s�Ol�Զ�/�m���{<��P��O��	q�H����;Us^^���+M[�R�?�_ӜN��V�;��m8����f��ַ�1�ϓ���~}*|r>�O:dZY�~Hܘ>>2͟��5G^��v��#9��Ϛ������'��$�Ԙ�,JG-�m�a�~�^�����2�݃e�as4gPL�5)�bҷu�*ޢ�m�����>CF�s�ξ�
N:�qQ�n5����-��`K�b�	�r(����	�Ҕ��t���"���7�&�7~#��a֎i��*SX%���� 5]d�F�9Z��v���D�?�9����Dx%�����gw��f�R��2`�\�О�B��Iǎ���H{wtE�7l��^@�n}�S���������LK^�ʝ��)����P����䙻��8m�F!%Y�����0����eՍ�U���\�?^���F�YQR�kK���q�A�H���d@g�z��z�H�h�h:1FI3G�+X����
t�h{6�b�F�����sw{t�+Xhd�v�Ш�}�p�+��UڥV�}��z�ۂ�o1���ʥ�B�{�U�4�G��95釸](1$��w�Ì<g�]��nI����b��f���f���p�mX���F$Ϳ`Sy�����t[�p�40dM���J�E"��Wz	E������\�o�Nə�g,>Sd:y)�(���VO�b~��{��Phx㘀�T=�v%\�fُ������͝�5)<�Ir��+薴����!]CP(􅺔�+ŉ�`*{oO4	(���]�P6́F������u.8�����F9��/zȀ��g����p5�l�&����pɪ�%��4d�>lUP���,�w��<�|��Gr��b@:���\�ݑ��Q*��}��@��ޙ�m��9�;
�<����\�k��W�<���iZ+�ʦF���cLI5=ފM��N��=�<�Uo
n�K~\�H|MQ���P'��x)�؞�QyC����,�ט����w�������c���<iJk8�X�K.�[q��O����*𽈎��JU��m�,9���˻�>�byY�0�N��	-�3�����|��cV,T4�{���n���Л�خU��Վx:�8��J�n���ZmM�g��V����|�~^�2��ꯊ�����W.�A"�aq��q"43�eq����}b��zk�Ǭ�߯�����A����Wwm�#�1u�N��>�㋓�y�k�_��|�[~�-�9p��'���mA������Kt�lE����)h����S��V�Z=�^7�Ӡ!S�������TŒl_x�24f�L��\}�� .�#'�%4�dI�/8���d��@|/Xu��gl]ڽ"���Ɖ���;��p���s��R-�J����&�缾�wS�
W��e6J�������=�w����hk�?S�*�k�]�Z2�pK������-�ul8����Ƌs���{��T�t]������o��Z�긚�'�����,�i
Ps�e�.b�doN�m��SZ5�d�O�0��%�!�>��eR�dlv����mB������M�qL�ܿ�,�7</���Лp�}�N���8�\,z~t���e��yߚ�4G6^�"�[�'�ָF n���hk
9͎R�~'�����Ŷ�u��%�������)M �����d��-�\jqS����T���+R6�&Yn��1����L�l�}l�
�l������ߘ��������>�.�o��Ã�}uxx
p�v{����`;���%qKZb�����e�@�;�R鶾�>n8 P�ʻ8�����D��m�//I�X �* q���o']�٥x�|���B�
 �H�ɗ���X�6����e}��]�3˰'��Ӗ��ΩBE8�F�_�(�M�ce�U9��#�����7�'S��ˏ(.|l|(c.ge�e�Pl:/�4�2���xb�K&]1ݥh���{%�����Em}Ո��}3�RlZp�J|*����Cii==�͡����zG�˔�����L��a^�;i�^�8zy�OO�.-�_]�>�[��~��̽��H�@���(��U��mԠ8.���~�g��-�;g�=�W���9�]�-��:j�h�I����m� #���c?��nK�\�N��<�'l4���ID������ܒ�b[��!�1}n�ٕ\��	8��n	�>���\��lo�,��A���E������� ڧ֖�^5��9�������OQ���}á�%����c3r�x�U�In���s[Qz�w0Y}q�碴Y�����/|4��������R،�h4�=@�a�n����U,�h�ۏ�����~[j����2x�F�Tvn�M�v��D{��"����DK�AC|8YYY���?�S���?�˞)¬�f�@`���^ 1����S�mlG$����)�>�(�F�W/�>
�[V%��@����h�s!��ᇯ��'�a$G,6�Q\Xh��aśhN���"adD$Q���N��3U޾UJZ��Z�,��R`{�V�^^N�@��������;;׬��abaFcac�.y'�h5�L���c���:bu�c�Mx�����~�IC;K�r[t9�J���(`��+�S��@��i���skc��Fv���}g�~�JD�u�%���'��F����.5-Ĳ�KLCy�u3[*�'	v�x"k'd��%Q�jӠ4�j��O�q��
f_�[f��D8d�?b�3u��\1�Qn���$�r��Fy�}w�i�(���8���y��D�'�\� �\���\J|�L		�g�T��:Y[��	u�A�����斖*�Uɡ1*����&�b��Oo��]:�,�����擲���L'H���EP�"�ot�5#=�����Ԩ�׎0�0$��dQ��ȓ��<W������x\ny�8l�&�hdv+����Dc�r�e�
��L:���5:����yyd���	�b�������q�<�A	A��o�G:�W�2�d4E^�7p�ʴ�nT������٥c;/����"��]54��ꁎ�/��/h\�%�s�����?�W?0�i�U���	�0��8Գ�34~Ƚ�� $f�?����c_��V\��Ǎ��N������ �f[�L����m�6)e�����]&گ ���-u�dK�.����_,������Y�칏�-������T�f~@�K�-���c��%x�f�!�e�<+C-�6Sc�u��)U��t9�t��4����[g7����\�Uh�]ͬ]����k�^�}o�gsqw�ki!�k !;�:���ׁmԄ�P����[��7�ayUUx��O�����&�zc�|����I��ǘ[}m'ݩ��6jt���^:V�4�T� ��0�3��ݧ�u�`��\�h����.MSkA�T" 
�)26��(R��ǈpC("-*�3h����ՙ��l�iqѴ�5.2����s>˷��X�#3��@#N�%I�dJD�+���� �U �>���Y5F�A�SaZ%�h�;D���0��Z�Q�K9u?�k(���ʨ�f��P}v��Q�	k�|�6�������#Z��ؗ�^_���0�����c�F��D�u���xzT�ً����$y�"���7����vU��MNjLaOB ������W�����h�ՙ5�E3�Q
'��v��"-�K�w�ĆS��(`D�'����W`Wm �:�H�,�;�``��Zo.���,K���\�di�d���r � ~�C�nB��nF�sss�l�$�P
8T�Ȟ�,�X���Ԅ��8�K6��Ⱦ6S4����Xu n~�O��rl~rl��?�"'':i�Q��l3�\9g~��+�:XX��0(=\�`�K�q���M�� ^�1}�Z\��
fӄ�P��S�B�.��=���U�8I֒n�r�ґYBo��N��=@e&���i�{.8�Dm��抰E<bF�(���=���䁋n;�Y��-��ba�τ�b�"�h`���w��Ld��֎�F�����-z��l�R�B��I��d�
�Pd���s�ZA!����p={(!���r����ZG �L�=�/�3�7��!!(,��h�J���{�B���ʯ�¤�	�Z/�΅��&O�+g	v��(�w|j*��vJ�@~���J�&�'���FO�n��R���i=�Ȃc���<�iŶ�r��E��� �(\S�R�].���|$�\�����Z�x`>�����E�n	��~�!�d4��|Ohu󇍡&�}�?K�Yf�`ۃR�����	�z�˼ܛu�I&�K�?^~��s�Y{��hmuZ]u�d��VV���C�H�Bn�`*4���¸�D��A� )d-�=��6Q���)<�YK���$��n�YuS����))�1Wg븑��c�L�_kve#�D�Wf�i�g5�p*�˓&j��R��X;.���	߫*[7${k�ٻ4�����2=&��m މ�o'+�&&�v��v�N�u.�qs���ꇣ]�V����0���e��=��b�5���VVLG�4�DsB!���2hUR���ӈ������542_l��������1��l��7�@���R�+�����ʸHܼ��/"����lmaxP�VbӨφ$��h2 c�Ud.��!�?�~�!���78��+KK����1'}�������Ss�S�p7��k`���`)�k�J�;h�(�j�G�x�e����e�X�P�����ѯb��@8��~�0��nBX�$�f���L����O:�m��8�r�$���c*/���o�\#��m�NJ��ֲ�
�������W�·��=Ӝ��1n,DRc2��� �������5d8Ӥ�I��O�вx�	~�!�f`��*�����(��B�P����J�QJr��`#)������|U�Ю����g_Q�*���0��H^{<F ��^��5��f�D,)Np��Ԡ�a����n��W���ë�G�N�P��qݒ�S#�[a-M�J�,��Q��<�v-�O��L1��yv�TXe;��
@-���$��n�*�@���0���`OP��(�/�%��}���F{e��7Y����kҗ�4h���d�8Q�7�����R�����Gc4�υ&ma�\���o�����q���\&X���
�'iӈC��:,,������"�{z�����L�+ƿg�݇�o��L!�~Ǝw����>�4���%ڏ�	-�Iǀ+oQ�˔��#���������&�ca�4y��t���;�?�W~�����?[��u�߹����*����)����̓[�wFp�ӿ��j��=�qT�I�E���k�Y^t%�T�-
�(2���+ݚ��+�f�C���Xx���,����vx�W��Ayzo��O� �%���چ���\����#&R���"�m܁�K;W����]}�9_j>�O���i����
�to�!�:T����IZp�_ǎ߆++6,8�}�;����=�����g�n�#i�}�4�"i!d��|=R���(0��'��TI-q�xؼ�0���Q�z�d.�+�|��c�H��T��!�"êj���#;���W��A^:���e��-��zΙ�	4��i�HII�-��N���8��mf�ˊ��f�xU�?�0z\!2�'�[	x/������{>}r勲6����t�r�{�EFEB�Ks�󬐨�~z� �z�Y�W�ŀ��m?1>nkkK0�J��[��;��Ǯv �Z[�&o�,1-G�5kd��ǋ�{�skn-�p�:O��f׽��m>O�2�~����N���l�=N�4^Aޫo���&	@T�qBP5��`�Oa��0�/Mv�9W���}��>�шh���>��F�!	!���������s�aBP�at̪��ls�e�O���2=�[z�7�T���q�N��Q{�� P�}n��bH$��n9M�ǔ�[L �ۻ;���������7G�/�z/��b�*�)���a݃�W�
��߼�	�O�>m��ue[�C���3���Y�����]\�m��x_0���r�ָ�5�I�,�)bK��0~]"�e�~��5��׿�Ѵf޳�ߋb� �AB����)¢a�W�|(		�]!���t��3�+7�U�!�� Y�.°����S���BjZ��(�7 ��v`Z���V�?I�w��'I��ֈ�=�/�v��K��Gb0�[4�F���t�p%N�kM=t�p̫��Z	\���A��E � >�
z�3����˴R�����&oA*�ccp�X�lw����CU�i
�\i��v��) �=�O��F��19�ϕj�\N��nM�Q��t��|���z��Z آ/�)N~`���J�{l�ɡ����畦�3s��?�|���.�A����-��4��X�Ҧ���v����3�J�a���EM���8���8I+�g��Y��^��N�C]�	���ThJp7�"�\:H��	�ѷ�WU�����w���!��(&&�d�Z��ٹ��˅(�H�܍	�Tcb�I���O
�l�aE�Q�*ue�t��_�X������:z�Zo��m����/�yB�o�I\J����!ʰJ��֒AjYD�����~	܏�`
���Uߐ�Bi�R�&|�6
�"�~׭ؠZ�[�ȧyu[�7��ء[˪� ��L7,S�)�!Lq�,hh�f<�*��.��� ��m6�p��#�D���n��Q9����H0��G��I]LZEZN��fD��8�͖���S�v#�in,�׼��c�@|��a�oĵ�.�kNjf��ΰ�v�А�����l�|^_���u�������ea/�|d_z�̮�*�chW�>���133���o����xc3l�
ņ������͘�e�Y�@��o�yf(��.W�����ʆ�m���j���/��.'p~��[�+��B��L��%�\3z�-�r~�(S���&M7E��[��|�B��?�3����,�����7G���^dN�/}c�3f��Z03���}��u�����v�q3x?��԰�Y�YY0���ͤj&J� ;�2֒�l�p
��Vvv�^vV�!f��)��.���@�<՞y�20 b7��$Z�ʹ��]r[r�[|�#���<�-F���҆�o^4n�Ko��u\��������6�&Y��D��j�J��l�ֶ|ww�֣�Az�*�?����M)<v��g�'��d�}����[D&�F>^^p]!@�o�Л��I�ߺ�� ���%�NK�;׬��E	! ܲWm���
�*����/ݍ" �)� ��"��Ҡ(H]����D��A���;/���1w�q_߻g���ٳg��5�T�g{݈�ϟ��:�Z(��jU�T���)��߂��WJA�0먉83'��'�Odv��u�~���-_V����Q��ܙ3U?�xy�[�
��k7�������!�5���f����Xy����I'E<�WW۽𶴆���G�A��1WWY9��gm�h�:t�����.�"hRFٿs�����ď�f����s�v��)gc�B~�5�eH/��p� �'œ���� z3^��
�h1';��;n=|K!�J���Z��ݧ�5����1�o�S�f��{Wҁ��	a�Q��6��p��m��HM�S]9%%��SV�c��Ʃ�#�h�����z��)�̬���X��q*.�<O�<��������
�a,�0�3�t_�[?�X_j֛��5�g�����K�k��qO44K��$��NE�П��-u�_�D!��[��$�'w��=F��;Ư�F���A�՘ ��	g�IZX�}{֕�ض�� Ha^��X1müX�z}����7s�X3�'O��0��t�^V2���T���MR�O4@�zA����i-�U2������_�9��v�z_s4���Z�^W�	a� ��,.�zJ�Ȼ�)xT��,�J#g(!� � 5��db�>@����, D9I�����O:[��.�n.j.�����*-�uRw��X��p$~��i��$�n����������t��i����	�����.�
Y{�Z~�`k������R�=#����� �ڭ��|�?�1�`����;}�d��St��̳Z$;��t��唜-�����]e:��Ч��ӓ�����[�P1��&�PE�f\Q�e~�l�H����3>�a]e�F$�|�Gq!�y���Ne��bD�j�8�l�$�hW#7:�Gm��Pބ���̵'L/t=�)��;g���>t�})�c�]��E�6"qCΫs�U��ϯ���ï�ő�Y-	�Ǐ>�),��p3����.���ֺ�/}+�!Ұp���B]��x=`	�f�e�	���B�i0��ˀU��9�6_0�v�fg����ؽ�2�VR�-�?�s���i���T��v�}�����Ϳ�B��``���D)�yA��<,_������M�Kꥎ�5�J���=��W�Ax����&�XyKA�qn�o����#��D��j��A�t�j�Yy��c����|��$i�ae�G�� �� ��� t�V~0é�1��tL�'z��H-�F��Uu���΍���~�aאˌ)�Z�+�=��w�ҡuv�qa�]�~ w�7����4�]��V��U�}�I(k�F�����}�uT� �D���=�����ā��^F�3�����8���[��E���Ʊ��tHt�O�~7
^M�!��� ����h�u!�h��P_��:nM�����v��E�W���H`xG�쩻hף�1z�����YYL��+$:X1�t�#+�!]4�g��}[h@��V�g	�h�-֏4�X��z��y��L�PU,!!��֙DPx��
 ���E�Ǻ����!�NNvwS,���?��P�X��-�ڕ~����є�� �[��qzͤ݁�����A@9M)i3�o+��.%%�K8����Bw���ȁdӂm-tJ�)��P]�ǀ��F���Y�	��_�)!G��\�a�-����9k$�zQP�I����@X�`,I�3�w�F<tz����bɨ�QS��Q�\j�ܼ��hR��n~#�p�	Ob�>Q��^��	;�S�0K�S䖎9r��X"!%�뿋��������Puk����`Dp�1�����m��F�4���,?��޻
S�w|�M�`�p�-De��b����%`�^^b`Q|[��O�3��{޹s�t��3�*��B8/����a������&�&rҪ�|M�.�{������,�GB�/���-��<�Ѫn9���5l� �gff���S-�8tj^�\�|��v�!��i�G��ܐ7a�����p�ef��L)�՗�$E�gϰ�u��mz�� '����SL1I0�M�G՟Ϭ#�����b����G^�$��uQn���fswFj�f`����lƉq\��1�Je�̸�]m�i����8�0�F(t����H�љM��1�5u��IW���#�{�fo�O����p���#��Wl���x�1T7�l{``�Ǵ��Bk��o�tf0�i.��`~  ��>h����6��*r��U}��QXXx:�"�]{�z�q�_��՞k�sa���2�����/����@�� !3�L��p{��f-+���D�Z<�]#��jr�y�驩�2/i�;LL�D;�57�/�m#�h�Sa�KHL�]֑�2w�/�� ����Z\��I�W�7ݰ�hӟ��~�*H���8�OɿA�hP_��k|����g,�N�)U�MI�ە��*ܛ96��/��B��d������%TU���W��uՅ��ST
aď�)aI4p
Y���v�߂��9Q�i�#�+6=�V�:`K�;a!�?׳ޗO��no[Ae����i�	�6����ĝ��&��������M_P�V\���n��yyy��}K����D�}�~�����P��{��^@#h�l&�������;廉�E�pݫ��`׮J-,�]�5'h1�(VI{�2�ూU��#f�3a���S}�Q�tl(mc�f���`MS"�>�~5�e=�@Ks���=����j���KQR�A�uW��4ך�R�n�{�=9$O�|soϋh}Ua�ޏlBe������99������#��4>Y���z�L�������%��)�eE����9�iшl$̒�'mW��|��̡tW���\�2�t��ns{Z^����٥��k���Oũ�{��\�Ə��L�h��r�?3Ĺc�Ԅ%/���`�F��= �4��r�x��t�H#�U�H7B;��̺=ڮY�(�=PM���L��>����Ђ^I���|�ߒ�a�3�A����ڵ@G�W���К��z�E��׵���;:K|��~i���d��E���b��ۭ���*S^}�Z0�������guRRXS'k.cc���8�z}� k�%����v(�ڍ2�d���&��m�e��P�R�vq[3�N��ԋ3�3!��8u5�É�6�4��n� z�}G�a֒��yc1_.nJ�V��C�o"�S���7f;�ӧ�\�5�4L	������A&g�~Ρ��*����Z�ٜ�Zu��+\4��b�Nc�F������ޙ�|�����R�1�3sԤ��1K�1E��+֊�����C�w.΄c,}G�9jJ��(qN�ւ`TUS[�u�i����T������[�#����0:�!(ck[�7��<cy�з�̯��N��qOO�徔��i�գ��K��$,�=	�����ә� �Gߣ�q2h��R�6�HÝ|�/�/�,�a w=���H�A���;m�|�#$K.æQB�����0��"��#�;�Շ�_~��I�h�R�|��̋>�"&Ts���'��̣@�F��\�[��a�[��冕Z����.�8͵��R	���:�6�J����frC8���P�~��Q��ɘӴ׹;L��>�b�s����feϗ袕$�����w�׼��x���Hf���ˉϷMJ%y�"'\�X2�^�B��
���{�Z	6t�A�>c�\�3W{���+r2�GnU�,##��6���f�;/QQYٲ�r^^8�6 �SSF���Z20�e�������}�L����'Q�ݙ���r�:�k���<�������-��~���JK3�ѭ����E^���GL�^���+k�$��i;��a� �Ԋ
8S��1�K~����n�%�+����[��s�-�]���d}�F?����hi����\YW7<4�I5�KLl��o�A3 �%��q_Y�P2K6��h�'Fk�l�{�dl��� &����秈�?l���mL��;�]?��2���4�J�Hܩ��A�cu�p���������I�Eo�+T�s�-���%���\}�cag�1�}$dt;*����V���)|4���˚��2�b��-޸�8$�c�b��<y�o��+��Q���B��F�k�w�m�<��T�O�>u���P��5�#''�����@�ʊ���@��p�Ǧ]�F�9Da0OGIG7�G�]�G�f���bDf���g@������5ϲ��[�4v�&?<	�Y<k��g(�u���MXF3et���W<����%�����>)|����Lã��]g�����T̰��8]�t�T��\�	%e�b�G��V��P�E�M�@ Jn�.a���w.�{�4'yS�AB������W�K�?�ؕ�R]ܾ�x��r���8HF�g����IX���g��W�N
��e^��)Q�lQr�����k��c��CS�6?ڴ���U�+B���E.je.R�M'9���^@�F1��l��`z
!��8�oLL��z8�V�qӆ��^��� ����CJJ�2���UV^�707	���+�������*���G�{����%44ځ1>ٞq�-�?>N���wQ�U��>~oX���Q���c�I��?������喝��I�QjԞ�B�0j�Ǐ`�8����K�t�ӊ�����~f�� �e������qK ����|��|r���?D��O��Th�[��b"ʔԬ���˽���y��L�d�wOr02���eB����3S�L]����Hj��˻:�����Ҍa��%���6�S�5p��X��D��ê�5�K��F욋��B�&��'g�S���J����'T�����{�Ԭ�b�)��o��
B��b{S5�2ql�gi),�Q-,���P��[Mr{������b���+yy>�ԑ��ߑ�W3cE!h������)A���eM�{�C��B�p	�A����^A��w96Y�Ⱦ87�k?�]w#4-*1]]�>�E|�JC���So~���{�^����Z= t��L��<�'���Y��ﴏϿի���(�\J����,�L�U�9������?T�K
)�C^�`M��Ϧ ;J(á����5?�r��yXo�7!d�!**T���%�'�LHv�Z�d�sՇ��Ž���3�C+OB���	4oL�����g����3��uW��̹���?Ny�z>�LO'��M~�.:xN�U�H�M�1�N��'�Z|�s�ovl��o�"�χ��$�%x-i-5#�f�'r�'�$�b��������o�����oGJRDB^��àr!`�SũV�'k��ЙŪ��3����x�4�Z�-X7���({��)�`+�`�Z���N��K��E�K��ǚ��(�*!5�e�D��xQy]m��c���䊖~<j�CG'x/|��E�����˴ՙު��!����G����5��O{����Ѵ
�>��~����%����s�.�����̃_i��jz���l�)Nc>����s_�F�NH �:4����+��P3230<�!`�!�Od(V�*W��oGݶ���(HeKJ����6ڟ�zV��&OJ���0���m��z�-.����g4���ǎ����i+�[ ���H��Қ�|(�Ց��.4V�:>.n>����5 ��H����y��l��	KYGG�0�ƻ�l��>���X|usSآf�QZ��_@@���3���p�Y�Ռ��~=��r����t�Ջpi��W)�a�N��ncsLa�"�p!���uH5�K>��z,��������C���,����M�s�����%�c:U�nB/~x��~_"Ǥ��N��h��+���ȠF���r�~�jH0$+���@q��YW,��{��*�lS�P[�K�g̊��PH�7�[�!������~7Կ��ύOB�,����*�������	4��v�JD��d���~`fF�[�Ck��r��y�$�ֵ:�����S[ɇv?��ao߽�NN���'�hUw�'�'�?;;���G�����F>�}7��hhh i��-[����	5�=�3 �F�6���>�#,,�9	���v�L��A���J�(����1g���F��:a5j��?�����(/��B�&����r!&J�
��y�wNJ<.�k������e�o�������h.U�uJ���wK�8,-8�?������	 W���MM���y��Ӭ�R�ڴ�۷o�'&\��̡ҵ�������CWLL̗zz����k.���Ձ���\	u��Ӄ#�>��M�G�{g}^�I�!������G����Ñ��S�y�z~q� ��ۑ��S��,�%���=_���1���fN]��kw!ܯCƨ޼�|v�F�-��o	���5�v/�_ݵ���V���)�ac�����5{N���a��m����v:�L{J5�Dw2|\ѧ�%�*��Ü��CThT�^ ���`��D1���U�1X�O���^U�|����f�[p�`�qd�P��xx)���T��>zU���K���h|��knβ��b ���\�ؐRT�-x�&Ku���/�ܥ��-���N��7H��I7[�h3����n�j4y6$��� ����`���m��r�ׯ��� ��S+	ߓ'�Ӱ�]'�8�<���@
�@>Q�_�A����G.����jU>Q⸥�ܠ�9^z�G��#�ѽz�
>�S�x �4�;?�������b�w{�n�U1}xN�V����	��a�K�;@�N���72��DB�8��G���d��%[��e�
�T���@�]]Ǧ�y��8 : Βn�����Ӹ`@x��GD�:'��GD@��:�����FFƚ��B{�MW8J�g��>���o0����1�]�_�᥊��c����lM`�N�
���Q����M^�w �O��"'(*++��QQ���M�Z�Գ�$?�=�z?a�I�ug;���I"?��3��r"����#Wh��G	`��y�����t=\���dddP��)^]9�y����_�9ƪyg���?K�m=����?�%�=��E��(_opV�3x��G�ϭW:�C�u<��|=��| ���z*���J>�ɛAH,�{LZ����eT�>[�����w��9�����B�°�y�t�[�4�������6E߂�YV�>r�sJߋfm�h��� �ST����B	���]NE�+�/�-%��^Wb���;0G������̌�R_�i����Xm.���j��ni?)	w;�c�����<G��pa�|N^����yI%%��+�	�,�%S[�VN�Ɛ���=�2r32��yB��Rϝ$T���f����aI�����eH$��j�:>z�]N��Bֶ%-OCغðУ�]��g]D��1}BBN5����}\|<�w�GiلeHJVV<	]��w� ~�VU����;��zs���|���,�<��Qutա��R�K�D���%�j/z��=��W/6�AE�oM�w�	b9 ��O'	)�4b����$��F�j�/�R3R�O��ÖԞ�f��v=w����\�M�uc�8��H��LHϴt4�/Rbo�쬞�DZ��N�O9��_(��$�t����N�5y�Gc+���e�'���҉�ЂBN��$)�p�\���`�x��m]Z,hck�=M*���m�a���3*%O~��1A���t����P,|�Y8��PF[�dYi��-�»�w �K|�g!�+3�A�%g8(D�FqS�8M��Z4������||�Ư怣�R�RTn�� o�5����MM}���X�y_�֟��^�-�H�锁�x?o'ۭU��������߿�Vd ק��ze��� Rκn�����>�U��[aҤ y�/�Qe���Ҩu焎�P��ǹ��L4�ė�'jpF�މ��x�M��q��h��tu�/v��s0w�� N��EP|=��S��SY���C��Q�-��||�E*���j��a��0��Hˍ6K�PIE�RRZ�G
P �972_&��ѡ!��9O�<��3w�$�/6ˡ���O�i"���������d��Lq#�\9��b(s ��+�� 3#���X:��7yrtl:@d*�72��P%>Y�s�c��!�n|�̸����4_#5��4�U�+��=Y��.M�g$�]Ao�4�&��_��0!�ƦC䚢�>.x���>P���9��D����Ϥa�;����ϳ����O=A*Ey�E�6��Q@JrtHߗ����4C®��Xg�W����}�m�w�5̫� /+�7d�0����KE~��_�wL���	 9JO/g?�����sW~
\�7o���[�����cs2��(�$�p~��K�?^.�ZקK%� �� X�2��
��S�z#
�ѓ3�����	��v��GO�M��Ձ���S�˛C�եS
}�97&���J�{5nR���W��W=��hW�bs�Omv.)WR��v��w���A�V����B\\6ߐOV���*���e���>��&h�;�����S�s6�i�вN��L!]S��@hj���'#W�Ѐ�r��q�?6�B�'���RF�ݠ&�e�ѭ���Ӕ���=���U��v�ٍ��qq ����ޡ��&��/���F{=,;�[[%�]V�N/W��R����]��7�g��TS�v��;s�c�TΚ���n��P8`yM^7�8'�������W'sr�h��J�?H�4a��eU��Ed0�(k�ZW0PQ��jDի�*�
s��:��-�9��2��5��}l�f�@�huk+i�I��u|��J��I��xER���T�JI�̎�F	1ƕZ���r�ʴ�ܡĮUi����G ���#i{V���>Fď�_��1�{���m�8]]�Uh���s�֛!&�����:��89���YB�~����x�ص@\��N�		h�NkQʘ����� |����8���OU�`��M���W�k�k��.� ,�U����ee1Y~ol�*��7���6��FKZ�P����բ0֏t��O�g�pT�����(�ƀ��.�	�ĪP+�)E��U<[��9��m��<�k���kg�1�q�vS^I�r-���3��DSP[QsSٞԨ����XF�#��)�y��G���Ma���ש�4����BG����%egg_��	�t����fE���*�C�� k��SS����or.�{�5�|���8���?q095e��Dk���x]�m����*P]]]�[Z~;>KOO���?��	��y�/J�C-��[�1g�󡶝8U�`��e'I�4E��(I��}]�.kЪ����Oq�c���������g���܄�,'|��%���2�3<�}#��a��R_���I�e�n��8]0܊���ö����4�F����!��tK\�0p�c�$���;�6{�VqRRR ��3p+��!��aV����7���x%�ܾ//T�֠��l9����������DI�ﾗ��P�h�D��U~0��	�CiN���>�Ϟ��7R�#�G�q�#(�
-@��6���%�_o�Xw��w#@#�ۭ#�� �&�ߜ��ӧ�8O9e(N\ӫ_l�l�{�I�JL�	
����>B)�{�ȟ%UB�Sttt�L�&x�%�G�w���X����^���Ĥ%���Hg?��V]B�^(�SB�"�u[�P�4(	_&��q��m���y�'�4�|�٨u=K(T���qk1�W�WTW����l�t����*�Y>Q �.�C�UH$##���${�ZXI���n���v xП�g���L�d�����D�r�MοVF����KW����fT:?m�0c%�wCy] �RYYY&*l�R���;�f���#1���̟�]�ޗƱ�h��-�|�{j��x'z�����2|�ݏ��Xh���-d��_�Bxe�(�p��L
8���������;��ܗ��C���fD����k�
4?C�K��Im��`������ ������>-Ï��f��#X��#��#Lp��_[�� �9ӢJ4��� %lQ-�MY����lmm�Y7�%�m[ �CH�P�'����p�\O��7�8��A����=J��vz=v�ڀ��Qn�\M)��';r�$�BY,��Y̴��c/�eM{u=��r*S���/w%�x��?����'�x7hK�n�>�2c:���������a�γ��%�ł{�V���(����GAW;�}��̛��)��?#��g$Q�Q�|n�n1`�~�z�P|ͽ�vR��,�%y���4dd�:�y�}f�D��x�_����ujE������ �ml��s(F3܃�]�H�'�U��Eb������@���ݷ�2<�������2�t���i`��7b��jj6�d �]hb��8?o��uT9�2�7k1���"�$ l��E���4��A�\ �^&���g��_3"���?NA��q�6q.��]R$l�Ψԁf���1�0{v��^��<�صC:���$��E����u$7,�DB*�ŕ�S-
V�)���q���\�*JJJs+����Ϧ5:��%a1�YO��m,S�*c	��8�G
�&'S��_T�����!$�H�L��q���%��	�N�GB����p)���O��̀S�^U�HH����v-j�VvW�w��V�-��N��q�����*���<��O�4�i����ލ���e6">Y���3>����,�_}�6��i=;�7��o���e��t͢'M�qy8�2�Kmq�ts�Q|+���,��o��]��9���������`E	��)S�������A���f8X��&i��w�Xo+Y88 a������2)t�	���iz�z"
h���J�8݋&NB���� �>��Ihkk�XY���s�zG�o�o؞e��n�G���p�$䴸�N0�w�9�<��A��������l�T'��)L	�I�*k�����T�h1�l~���|�E7��ۭ��vE�kb��x���Nݦ-`���(�\Z����ص�Z�"*<͇�J%Q��لݗe߇B��a���Y�>44)B$6��0|\G.�0�R;ne�}i杚.(]���"z��Nf��5]r!�Bۢ�.�:��z u(����5�K��w^y��mU��N6�no{6Q�.�455���	_>��[���N��
U��4ݡ��ݠ���[r?�W�w�HGO�P6��~����X�n2Y��.뗗���T���a�.A�w0�CT��o��ıoQ�����e=�0x�����L��G�P�
Oۖ1�m��� 
:�A��EB� )D��0��ChBƱ���}?鿿o�#����6V��{�i�@0���_cY&� YH�"�������B=r(���;)����/�L�gb�zY7�� ���@�=�(N��D��d	Yل-�能=O��f��DW��_
0�Nǭɀ�m��s�W�,��,/M��ܙ_�B�����JV���1%�d�K����NNN�Bs�)�j�MTFR��ߣy����UWΣ"H�+���=�Mj�W�Qiؕ���|}���)-��ʂWՠ.���^�F��i�]�H�;	�3nkg�� 5b��EH�A�\��V�K?��H۵�H��v�~��q��?R��O��ښO�A��׹�����CUi�8�
�Λ��4����t�tCɛ������r)i���L��H�{�� o�|\q��?���~R��鋤��1������ mP/�H�T"��- G?5.g����q/෬��o � �7�!���%`�?�|�ص ;09�h����0�r�4-ㇶ\�M��IRz���Wl��I�?o�p�k�Cϗ�ME5��K�6��%��}�'??ߦ���ْ��"\�2 ��ޝ��&���t>]�ߦ)b������	���8w�]!*�@��Z�E)Z�equjG��0c>Z��%�C#��O£����B;Һ�3�{P�V�Jr[JU5́o�_�=�����Z��Tl�Eڃ'���*q�"+��pqe�{�F6z��{�Ώ6lk�����=�Q�����k����Vb�MǕ�A��̣e��E��M��2��W�,h�A�Wz���"o��������r����r19�R���
#�#��F�$���)4��vb��wE��1-G��*"*%g;�$Š����¯�Y����MW[:�ܨ�>�Z��9;m׮,f%Z�tq ��0y�:�ˋ}�����y��O��ƉaRT{֋��I��To�o�V/٧9�nF|����;����B�8�����x882	�����v([|Ѡ� c=QĽ��'�CK:���i�9?%�y廯�$�D�7%l��W��l�JH���|��J��8�	��@��x�C�;�<�>l��H�,-�^�k&j�����s0ʷ>���/���9���eb��U�(4�쥈o��a}+m}b����K�0�t��쭈ݐ�"�3�+,�sq���@v)����ާԠ;c�:��d��4H3}�D�Py�K~���ǒ �%j@�FR9�oN���7�F���COA�&�˗���n�~Q���ݘggg�mi��0+�zL4�,I������T�6��ۻ�U�[4�"k�/lY<�^��Yu_����hQX�SS �xr���%���%�D�F�mPJ�-Y}y�e�o�p����)�P<c�	Vub�ٴm{NQ�uA�)�;�-!8�@�8:��p�$��%6�R��A�~�����4a�"�p%�=�KO1�[�_^�ʃ�j�����9̞ˑ�䃽Nj㡬 �B��o����Es��v���,�$�������<|ͨ���r�Ho7>���3�Ϧ_z�st���ix�����Bs~q�	�S����5q+���3I�?��.��N�8�F#��Y>�v�.���ܗ�Ӣ�/��R�����1�E��Z �'�
�{T%���_���g� �U��w^��` � A�-Qd���1��/^VV6�L�TE�>��!��Nyp����c~~����;�>}z�*/-�sbf�S��$#�f/c����h�#��y׀�5�d	dt���7�����"���!X����.W�m�M�,�:�S�tg�z{:eȒa�{�=�^�v���2��Jwm��0�����X}�BA4��b"�F!�-�İx�
͇Vڳ��h$7X�Z�H��$����	
_�n)А��iEii�������fO>�����A�2B���kH�22 ж���8!��2�^(/�����5؈��<���r��z�\!&�]����<�*N�@5L5���[ �}�,�o�p�ma�p�糿�mDy/2���!�4����h'��k�����M��Ԧ�����!cQ�L���O|�$F;�1��"��Ux�Ɩv�B�c�@!�ЁZ����q���CY����s�Y�Cj9���Él:(�O��ѾM��e��&�������#���#��b���_���E�^��i_A)���.R�o��eNi�Pt�G<�aۖ��&+�XX���������^3) �L4_�)�)���#yj����!PDh؜�y!����>����Iv�R�Y���������g7w}Ij���[�=j�K�$%%e�E0�,�f=��:���񢍇"���w�Q��X}iXj�oj��NXL7� ;��X�p��f��k��7=���]�v(>��Y�Z���%������G��߭���Sp"	���ug5,�W��?m5�h�;C]d���<���ք4����|j~�^�5
<�qV
@�p�\#jIn�#/�o�H�cf0ڛC2��� Z�ߓ�	����U0���_�G�y��O��|��;�'nН�� ���6#bB�2�>�3���X>fw�]1tGV�)阮�h�f��Lh7W�vN���J������7�bUU����PQ������3����]�¯�=����ɩ�iN�����ᖌ_=w��ώz�"x�s�|H�VK���,>lły[�:>>��y4�����@�Aw��2��*�4��Iw��<̂��]=�,�9��{	�Y�w��{F.ݟ�4����`2qz�8���03������ʶ$X�b	z��:9R�_z@0�:!���������J��ŉ�j(	뺩�R̝s�C	|e)�h�~��pR(��İO�|���Y[[�΅��{�	��4�`t�����*�(�AU#*�K�n��������@����%��uP�|6�.��pVm)�ՠ��t�(x���h�\O3IĐ�e(9��C�L�ٳ����zL4��7��2I�l]E�嘛������y�|�.��\��A`�;�'g?n�����&�_����I�S$�̘������H�?j>��ʧ��HJJ2\=�g�a
Y搈��ʍ�MmS^7�J�����\���1o�"a�#y}�_�	2�_6�/#����E�[�?�.� V�����[I��`	eaa�p����ϛ����m�[�y�!��x|Z� 5���9[�X��:�,�?���3٠)��u�N�Z��\�T����2b A�����#���O���",�ۯ}�"�囤ǈY�jϏa�-�����͑<BQ�+m��O�	����9�#��2��Z���Ge��RC��Ň��O�	a��P�hG����vM''>��5GU�@��4�=qorZ�}������F�Gng��9N(��x������^���ǭIJ`��g�T1���[x ��t�R]8�"^<���n����w��Z����32���
���,|}�U�99BoǠ�.Cu_�kA#�IU�����qG,u����Wz�j�>&���*n�>?��s?�'3NK�^�K�R�tlӻ@��GH.=Е�I�&e�*-K��vz�=$�W�LO�M��WWb�y���b�-�)̈�B�=//Z?������I�m�$��` xi�P�oKvdm��t���	��qFH8�Uhݑ^и�Q��>����-��L%2�ĳp��´��N��]׆��⠹���b9�N���/��W;^�"n��I�Q�"BD��5�@'u^�* E�c^��ί&�É����h�z4l��m"��B����x��\JA�5�78XV�Vs���!�(�� $]j�NN:}Z%N������#�@�)'�����K+��|ݙ�����$x����������H�͜�}��oi����i�>�>R�����1���z?�(�>}Z��"�]]��뭭[D��L����@N���`��;�(������y�Ɔ�\+��.��2/v�T��BѤ�zT�O���fW�ݬ9fㄵ��v���0�D��3����qd�<P�o�݂U���L(�ʔ��*c�Ujg�z���v>$3�}30>��<4��O|Τ��9G�{DUU�`k�� �U|����p]]]åc��qi�n?ړ�8�[��qk�g$7��(��o��j1���>E\�ɿ	w����F2j�4�����m��3�
|�ۀ��"$��UҜ�|�HN�G;1��]�Md�����r냗��quS�������A�����?�z�/�W��5f@�ˁt'�x���t��"�0^�Ǳ&LGGG��ot�9������gr0�5�5;${�!�t9�˰)�&9�0�\%a42?»�w[;.no�D���ɹ�@GX�����ι�vk@��B��F5'08�ő�V����u�۲� ���B���PVx�[JY�?�s��'Wb�1�S�y'�e:96��ը��Ą��fƬ<��Y+��(&1t���]���CE���v���C�U(����ȝ跸o\��7�\����-/]�m��F����,�e���r�hp�Q�Д���;�e���}QN^?��5�@8�L�@gNȱ�}���l��eu+�2ʰ���{��.������n8 ��88-+��I���Όv�l�+9Е�ʖ��$��<� �d��0�$ۖ��c�S������h�[�y�H�vY9�S@�����N����k)�u011�fB��7�}�n���-b�zq@�z�d�k�~�^X�߆��{���3���H������%Y��]��F��[�K���fq�������%�KP2���E\����e1�f|+�E��Z���j���P��-�ׅ�������hDD(�I�1��@��a�3Zl�K����hd��-}F��'>���"f��(2j#�L�&�50�������œ�_�GHGY.�C~��}_���h�8,�+���N����^�#��P�YZ#��,�д�R�3�v�X{�N�q�?��:����^RS
�;r%����o��wN������h�M����7��_;ȗq�^��j�V����mya�`a���!C����Vj&@�fJ��\\\�O�˦�Cc� ��-��{vo�+��~w*�K9 ��v�۟��(�W���%��.�O%�dY����50@��C��E&�qq&!�A��=��gԮ�y[�8��AFQ�]�����	U�����60m�k(|4�b�G�����A�A<��r�X�/�j^�1��IH'^�C�O�z?c�,c�^"��cMF��,�j��)lQ��z?@�b|s}�a�͎T�� �m�)g8Lb�,���n��:vr�(�}�{����ô�,��G�"\\\�	O��
������L[��'� yi�K�A��@�?���6g�%b�x
��vw�m��\�㋧��bL���ݾ����8���0�	�ݽ�t�賷�3K���-88�#PeKFCC���A�Y��k���r5`sW2r��!%%�Z�����3u�Z�D|��w01[�^���}���v�NU��s�g��x�#T�;=��x��Atuue��58:�I�]=�H.
�-�W�E5u1�Kn�S�d����I���}���9���k���[�P�ޤ��>��t���ߕ���⿚���gb/v]�a��b��yh1`P�Y�^ ��T��ⶈ�-����ϊ�K��oZ�=�aZ��L��^V�e�Dz�/..ʷm	 ��j��m+�J�.Z���]_��+ t���Zz�|��ML^�y�|os�3�����,w��승��e���o���z�#����E�b|Ǆ�������Q�XG�`�7f��Wh�ubY���	X�3�4��;�O���g��pH5و�-�r�b�`����Ս��vR����>H����N�A8}_�aT�L>�'��SS�]Q��a����)�!4�VY!����y���!���ܴaY���]��Nn]]�ZF�fЗ,������7�]>Q`�	�<D�+;}~�İ�P(���N%y�5 �n'�@����d��})�x�]7
kNf�J?�5�^׾�~�Gמ�����9�x�S��T��o�]�l���d|w�^�$��*|&fy��tϞvQ~��1�PQm�ߣ^E�t��tHK��tw��t34("�)0�t� -94�1H����^���b����y�{�s�y}2�Z�ms�^0w4AHL�QUE���՚Wwl���P^^~�H-�r	�:D�R�@��|%N��� *�C���mS�����A�� ,�w��c2m�g�����N7o������ò���,�X����- �km8�y]�k�������gO�hi�#`[\���"b�7h럳y퍾��黗����-���+]]�]��m��M���{�j�����C�}+[��SY�Ι��Ϝ���?Zc,�y{X���޾x�S�Ë
�h�9U�n]��A�>�DVYYh�,��:w��=%���߿�G�0�@rlb��Ϳ�����5 gNc���������B�s�{{���(Y�����C1���!�9�A ��ɉK����^�5�Jo��#SS͓�o�i����P�1sy/+/���!bz�k�؊�/ݽ�}���+�Fl��:Ek@*���� J�}�*��$�mU��K{'��cQ�֢���P���.���&�i_�� �_g�4S
�X����8�����p�{6�^D�N�1<,,������T9�o�z��r����(����<���$���RUK�ᡡw��$��`C�J3�)��cJ�	H	ş6������f���'�H+���ΐ^^��rnT9�����".>����uyhwy#��5�'�[������E����_[X|���{�Uo�����b<��%�ՙ��O����:�i?>^�M3eѭ�!b}�P¾����nn�Y��L{���"�GR��4.�M���⟒�ƽ�IL7�n�EQ6,��UD���Zj��t���-����6==�ck���{P�۾��9Q;nF�	�l�k�P�qXO�N����TM�>0�:��Qu��!�����E�L�-����V�2���/�k>,�3�$�H�Y�����~���5/��ޞzn�{^<*����K���č�T_��s���b��5vx&hY�>B�t�+.�|q�V��M�vf����;�/�У�*�f¶&+iXYoC�\�����W�`�>�>�j�ƠH����L�i[]Rj�`�h��/Dd�G���'{�!���jñk�^�ץ�ͪ����;MF�.���i�RDf[*��(1�9�y��5)YY�������w�c�0G���`�۪�JRű�4�di_�t�	�c�&�֍���ަϦ_�2���X-c�ڵ��B�[�����}H��?0?"d#{���<��t���5�l��e:Il+�X��bt?��ܨ���^��Ds�L������)^W�c�_'���w���ձ�����m���J�û�%[:����+��'��̳���c�j�O}}E+lQ
t+��8��{��ʐJ��q�څ"�3��Уe/0gs{=���Vo�AbzM���'�A�7�����a^އ��R5ؠ�c��+���}��Y܅@�Ԕ^YEŋ�gK��!	�A ����nQ�n�xi|��8FT��F�_7	��L8��c��J��/x�}�d6�]&q�ٿU�|�u��U�@��b�M��BBcbbn���`����ҧgV8�(|�{��_�������>�.��Շ�����GBz{��j*O��F/�]�	�����������wo���ߡ�ލ��`O�DebbY
����*ъ������{s@��u�w�+�����;�僟��?Re���	^�q�q�|����e]���|��[���~,��IE��0���E�]S,���=22%MM���S�8�L[s[Ҋ�_(����.�����J���I����l��O�b�AmI()%TU�ǣX�@{ʐB�~�����z,229�7�u(��~�0(�le~&2侥p��!���5�k*/�$+�o*"?"���]!�	���WRQy�������@����?�L������z P��*r�Yŝ���T`0��m���bq�����̎�:���~q1�@+3�5������'�i���@�*')D�Bw����
J���n�m�����-�Px�py|�X�\d�;]!�$x���'C?�����b�p��5f2�D�b"�#�tX��]����e|�b�����pZ�f�(���T������0���3L�g�]�����a����ar�����Y�x�3Ӣ��ܰ�_O���qG��mZZ���p2�cE��U�U���Ó�r���	C_x�P�=RH��&6�R~��i�Y�:��ۯ�A$��~�9P,)H����L��k���]I��^��'5�	=�������X D6�x��s�Ҟ%��D:�ë)B��$$$�/T��-F��#�L�4R�!����Ѽ�������|5�)��}����1S�K��h>�/��H�����:d|��f�b>83�x�����̬��F:4��� ��P��Ʀ�� ���۫пTWk�џ��"��!2��t{�Q��J�b����?�9=�j��p�-��6KO�b��):�[��>z����N�	�Q���)?^1ʔ���XGd�KRWQy(�)���g�a`�ê�EnW��(r��*}F2)�`f1U0�4 �Px�i��[6�3m/��K��� t?�>Ya��E|��qq`�MMLXY�)���
��o���J�_�;iJR��ϋ��@h뛛jpxeMm���t!��iQ]]]uC�"��Ng��?8�rf�7�����unO�zɮ�WM�2��=��^"�N!�bd�|����k5��d�<�
I�6�IG��R�?��{�}]_��;Z���c5.V�
X�(D�����?��σ��l):�2�&T=ڪ� B��:!͈��щ�i�f���ɂ�\&W��^����{�]K��t0#��/2N��}�V�L||��r_��əut��
>S��n�1R@Df��%�0hV�1�?π���P�vS`����I�����3�Dyee��W�u3�܏|��f��[��Z�܀ݻۡЩ�D��z��icfb�Ty��q��9?~)�ٽq`���P��uī�_�|7�lϫ���q륳Z�9)���ۈP��3���o%m���h�iqj3R��Άݵ ���� |�����$+@��g8�Q���U�\����c��Qwy���Ht�{}�6H����=�Тmt��n{ز�P(�.�����	����\Κ/x�W����}��|���S�U/w�,��n5�Â�<2g�RI�w� ��ڢ��Q�����,����S���8��Xuʠ^�u�R16� �P�3o=Q��=rM;y�����%�s�s^h���h۞bim��\i��.;XP9�+B����%$$�^�����R�F�����bx������Q�� ��>����Us7��g�=���Ū�k
�D�����1.�'�Jj�SO�����y%�tU2j�;t9�t1FT��y��,���50��
Li�_����*�N�\dOT�V�U����Qt,7�7_d�󩇷����̶:;ܒ^�_��355�̼��������Q�����z�B"�����`xw�j�����8����쬈>E���.A�5����-:::��_��M�lUL���L��dq���	� �4u����N���>��� ��,��2 �QN}§E���!�Wa0�w$ab���V��=��L3����պ(��!}O�t2��|�B�z/�K�C�L����e�a�R��>-��3vm��Ѿ2{e���nO.��SR�r��!O�A�����bG�KQ>��2�x^�x<j���p&�,�n|�%v��5��~������1�7`�[0V0�d��?���������p�ә�m_g��$���A��q}�O�!��JJ�G=�{���F��0�tv�|u����E�g�k=|3e�t0�{��ޏ��N��x��/j��'�t0��'����EF��2>�%�3"���,�����$,�FX�7���JlW�����C��kF&iPV���ѽ��ֺ��Tac�}}o倴('G�ǧ!��i���#  ���V�o)�>�.�8N	 ��v)^")��8��ibAC@��	�E�;�a��O����q.��v�Aäʒe�sJ�d	���%���\�?�����8xr�.�]������B�3��p��j��{��-(Pם����ܗ��8X�L�m���C����Fn�֎�f\]�Eտ�Ю�����D�7�:�(�v=v�d�F~uS�~�_�A���#��uk��1M��L�n�:����u��c���[���܁$=
��;/[�c�n���a9Zk�iu>?v���yd�B�f[��4r�����OH(Z�Z�0s����w-/m�K��T��fi��g��B���k-��j����� 3���h=�VB�w�d$�П��/'^�M�IMY�ܛ����A ���y��+w`�!������1��|v^�l-��X�|ζN��Rٽ�d?��[���8"ǧ���<cI�O.�8hZʾ�O�����������8�S�?q2KI��x����fPV]C#(�������8�㜳+����t�e�v��K3J
���̽�~��4���4�IP����*I,�<��~�t5з�BT6�����=���@���V����Z��ޓ�1�ꇋ|�y_��j\��#���a��È~`"+l���$--=�{�ʽޠ@��y1����g�pD����?Ж�vSqʙ�V"�����>[B3*Η[Z�ǳĞ�0_."�ˏZ��HCӲN�Ҽ�@<��B�B�eD06:��lZ&��Hx�ǽ��
.3���aԢ�	�5� U��!1fă=��AR��E�S'�d�`j�����F���{p�����~��f��s��M��mo�m }�f_�߳ �Zk*/J�b�ު����?گ��[�S�����dt�K��r<��5�`�&IRRr�jtC��˴�N�Ѿ��~����v���~�}U�E䨺�s�H�xS�a��T�ZU^�
_x)tӻ��|T%éԹ��'U����+5q�$0�}o�b8W���E����x�S6$B=CV���L^�-��خt�:��\\\������+�i�2�HB���zD5�� ���֮��8c����%A�B�b��T"׈�q��UQh�c3ei�ങ�.0��r344�^w&����u���[-C?j�I�,���h����l�4�?�SQ_m^�K2Q�:�=����{��e�qT���,�_�S��l�:_��V�����(+ۺ>L�r#��b��(7W���jp���9�Cv�(zőhM8���!x7�M��`c��(� �[cq"��	�����[9p�/�R4A�Z��>�`cc/��`��%áU���Rpd�<��@��t�ϟr!� �¾]��槑|��5R����|�Y��3"�e[i����"r�yTJJ�z�������N���B`0�us,����g!��Mj��u<����̬����ю���d��OK+��AY���qk��`z�A\�W�9{N�����ard�i-��Vt8��n�N� {�xgAZ_PXX�˼7�s5:""M��^�v�s��KT�!.��s��}Qh=m����Eej	��-�2h��*�����:�ؕ� ��։Rs��-�,Mw	`�5�����F�b��9ԫ,y��Q��^}L��ᑑ��%.NNn�Sg���!��k���3u@5����K��4�󊺎�/,�̚b��QZ���^��;��D���oř'��Z�JUSU� s��ꏃ{M����A�ĕLp��5�M \�£Pb!�]?#���:�I�B6dע�5�l+A�������N�=#,¼��A?�U66�1�k����ׯ^����4F�t�0s�U�k�Si�TgPtq�w95��R%�*7�K��`�r�|m��`�o�*�Ǻ��4�@�� ��L��2�ܧ�a���B�Z�v"�S?Dϒ�T����_q���ZT�y�È��yy��3w����'�z0:�wO
�ԥhͲ�A��4ӟp��;���*]�׳PY��ny3j �A�DR=����2���b�V�ά�<M�e{zz�Q�"�� �.�=��	e���������y���DII	��e������xl��:�.vN�ݡ֐�9�T�Z�����r�=��ֻ,�_�f[=F[?������\K!v@d���A�/6ӝ2���,�N��H�wF����q0��Œ7C�ڴ��_P��=+�#B� ��u��Om+'A>���<v;金H�����>��|NN���p������D��X�O�<���◵>�g�P�{��Keoܓ,������ �����2�����gĒ�D�r=�y���t��f�[�ow�u �c(Һ࠮�~�u���y�=���hy٬�x>�>ܸ���Xj^Q���7R��R�(�{�vD�I���nQZL�X[1D�9�6���CJQQS[�T_�#xY�j��U�*��ط�MI8���vf�e���A�w�T���55:R�&��<�S�!��l��p^U�^ I���;B��{֠��]�'
�|��-�rt��"c��(�����I%���YY�No0/�Zit�1D!��zL~_�����[SuY\��~��o�㿠�y~�r[]_]URUU�v{����jXd�-J ����3d���üx�vi���ޏ��x/�^���Cft��}(d�����~3;�������ؖkO��'O��dD����K��9.Ɍo����᮹o�텹����&rY�=�]�5�R1��/	5]�ښ(/�����ߤ�;�tut|� �����؜��}FϪJKU=7(�Si�x �@2���C/�rS�}�vUs>\����ƕ,E
y���5�6�wȜ)����&�Y@h�yX�`.�D5�jj�����K��u�z�$����N�}���s� �0�M?wbbbz4Y9T���p�ָ5Yy4~�������Z9����65��VM��M��ܗ��l��SDX��+6��Z_=�/��ս$#��4k�^� vP����Q0�@iD��n��k�QT��H��ά��fo</��9��Kr;jٕ��v�Sm��A�4\�=�$4
c܄66�78���^���;[�~�J����\+1��2:g�ZE�l�,�� b�~ v��q�W��\Ӑ��&�O���2�'���5�F��Exb��E�Dk^�D{/7�}R8��i�ˬ�+���G�r_J����|�
��_C���G�h��(���Uy���K�%=W���A���P�[��:	��rtttL���6";n�p��5=���-��x������Q�=EB΄�5�c�2�,\`h���V|�D
��`�[񌞤d��C�I�@���@B��:n'J�	�*~��7'#ø�x��p�]mCԟ���>ꋤ(§� ���<���} {be �K�,����ͥ��O��.K.. ɏ?�$����B�x��v��})�{UZf�=����F__��):ķoJPw�nȯՐ$u�_��}��^�.Lx����#jY���U� Q�w[KA!L�*< Hs�����\}��V�h�H���3 ��%G�DH�7٧7Q�4�)3 #NI�K�FU�^	  h�nk{P�� �K�U��SPg��TPh*��g������٦5F��q4��+)��X��+>�H�prR��yfhiiY��t;0J/^����6b�j3��H���[c�'�T�Sa�ڌ�n����F2,SY;�՛�������c��G�EbAx�������E��G�	�����n�k�R�ɶ���]���;����%�W�-�ٽk� �rۿ�CFc_l)�N�c�����VJ ��|���<�8��x��X rCc��0˂IXUr���x��]�;rM}m%%�<�����i���� ��F p������Gp�4�q�����qk^��FQ4�`�9��c�t����eW�)��\���4�=��������^;��-J2��:{{G$��3�8-k�,N#��>G���.��Q�;BiM�����+Ip&��}4�5I 0,
�a�ĵ�mw�j�N�ҵVb�! �S잩���7�[��-����-d1Y��Æ�wRt�
}��D����C�QZ����~7��%��z��u�GR�j=07�zB��i�	���	��6�@{�S0�+������S
�gׁ���t�+��� ��z�����݄�ֆzѠ��j!t ��J�a/���VZ�L��o`�7�8���y�v���[A&>q�6�����v���٣3�CkDg���N&"2���aecA�d8��^�S�ˌٷ�����-�@|��0T{������`W2
t+m������j� Z����${o#��}��ؗ�YH��#G���������K����(�S̷�v�Y_2k㌝EL�#��K�z�O��#_���q��s3"���=��Q%$$��K�[+#rbl�v!���?Œ�Z��� cRR�z�R_��XbN�\�쬬TMM���h��R~C�*�'�����#�T���wD/r�C;���-�$C���LC#����T'WAWn��/u7hե�%::���켭�.�#M������Z�����Ɨ�>==>�8<t������5��,���-u�hE���M�iM���_��c^� 1��UK��v���9iii3^ �+�fD�b��u���F߯�X:�O�)����		y ����"��[!��}ް�4m{�ڤ�+��եK똾���o�n}o��p�f�rFH@���AZ 8 ��0�����WN9���6l�w�^G�e����o\��5�I�9>�S��8L�j�(��%#'g��Ǒҗ��K�s[D�7�h4O:���|+��|�Mӓ�n�R0M �V����7:�S��}�i$F�ݻ�����hsH�RO�7j�)HN���NJѴrf���
�tI��VE'�K���:�[{%�*�6	�@�#��\����tx�v����ABX�+ /� �Xn�������W��MWw7y��́���K����S�:U�i>|�2��q�vY��d �	J�١�8Q{�cg��<�^�w�`
vP"\,�\[8>���90��rn�j5��?�B�A�5'�	��VOy6쳽A�t)��K��Hŵ���ƍk�ӌ��,���?�� �G���$u���|���		�	=f.��9�U���dCkKk�lfaaaF+pi�f��O�nYO�XK)3�K~�����X��`�]�
�ݿ������N���)��vϫ��L �y�K�T�f �f1RVMI�������۫����Ѫ�/�$Z���ā�j�ۓ���(6���QI�~�۲��)l5�BHDԵ�Ki�8���q:5�2!��
�9Fn}�������Oe���{�򤴷����oa�0�M���4HĻ�D�,��J�EdgK��Q"o�M�@�6ۺ���q���=$��~�PLK����n<.F�"7��~=�5V,rF5@,0�e��茢g&�F i�%�h}h�`¯���$�L$����i���O�����g��q�pV��FY�������F�G��'l>�s��	d�ff���7a���� ������6b\�/��:) ����A�.窥ބtt��-~̒�Jl.ϖ��jq���p�)aI��ǔBnJ�L���(�]Qu���76]Ӑ�����n����0�1��5�8Ӧ�Y`��D������ţ3S����'x=_�A��BTԿ���:bV%ElF]�s#�j�5z��Hi���ϯ+��0^tI��Q		V6��2j���>�r`����m5��t*�A|?���<W�㓬Ivs�b��p�����]��)vrV2�<��u>����9����,yU��3��j�oo7M�P��
 ���5����tx�� 
�ܽ���Y���8�yu����W IݡFsQ�Yڷ^��,���3�����(d^ƕ���L�s d}s�3-��9{�Dl�'&H��!A� KOn[�:�<���2z�`D�y!G�.�ͧ�M���P�'<Y�W���Yz��ḣ"O�2�Q6@���*�,���j�m5
}e�a��􁜇R�3��Zvw��d[[5v���8n��&(*�i�ϗ��>����-(����=�Ȯ=��?+ʝ)�z��/�U�.���O0>�����������@���: 2�9dѣ�s���������>�h��s�Ky�+/&>�����}~|V��{.�Є���S��u-:�S��]7!IRe�p �>R�X�3'}�%<�m\�9���H*#UV�o+�����Ԣ
+*x����p��}/={� ;��A�\ �>��F�2�H�����/�?��׊"�I"i��R_Hb�7�'�ܻ�ڝ�p�#4J����N�cWggg�	{����e���������"Fۿ�aMW]k��F򕽽���AM^���a�{�R:�Ž�	b�Dh�IIyϊ4؅Od����X�qa��
�˃1�!Jx�����D�iP�*�"�C_��*oMU���ʦ��7�����S�!��r��$�@�A��U-����Tp}0�OcS+j��ؾ��K�����-��b�o��I�"{�}�f�;��4�H�:�ѭ���*q�G�H�9�(�8;g�?�������u+��A�o�aݟ��[�W|XF���_K�t>S�$�Q]kC��j�<�l0��~ ��;�Jߣ�T�o-�;C����� ���M&|^�����3E�!_L_����Ȭ��޵��3����� �	�F%���{�Û�t�q!���3c���*������TZ:��br>0��*$���'�5Y���~���B�$�YY��P`3i�^vE�Idu[�D��#5r��k٩bX��x艉�Wآr��c���xЫ��	 q�+��WZ�Կ m�Qy>�j���y$�&�c����i�����cia���ނ�����GAZh�=���_c��ۍ�Е��7�/Z�:�D�yc���I���E5�bW���Q����	=s5"Y�D������JVV��.�� .�0F��,��Lq� ����Q�B�F�"0�����S����7Pl�b-9`$u����^7O�uM​|��6.d�!�֮ϡ�&{!3�[*}y����N���5w.`��2i����d� ��3�Ʉ���lR�[o��H�h���0ųw�{�	B��_P "Ƅ�,%�`�,�<J���S��4P4��xI(��7��M8���:зu�2E���_�Շ%��B9�#E�#H~�k�d}��m3^"�N��"�7���v����cK���)��hI�0���u'���y�eHT�<�k�����s�@�3H;֢���JD��6X�9P�1��������Yr���T�!�ا��HP��0pX���^fg���D�o�&x���}�!�0���n:��Nni)W�4������S�w�9���2TVN۾\�>=ASU۝��$x���&(0M�4��my�8~��,��	O�(=}��8�/�5��`�����T���dh{8�#P)�.�Ϟ�>�b�60[��9%}�7^ة���f�wk�^t���o�ɭ����_xm&2�@ ���YH���T�u_*k3�c6{�"� N��9�ū�/��)L�yX]Q^��/H����)J�Q�m��d�l$4���B�o�0�����v@��X���Tl\⟝<b�|�:X� XvᛂTǡG��9�/���>J��N2QY;c��ۇF��r��մ�)H�����t���0t���Z�hYG�2�&$+���M��
�Š̑���,�zyX0�W@蔘@��
��К�j��A� � W@z�["�Z�T��ߣ=�q����{�	ч�{���{���4�7Q%*�b�IxA4�"�FF4�s�iiϊ�����rsk�}��zUL�s�IWYjV}�����$��vǰF��)��g�(�-��_��i�	-AC
�p�z�=���S�s�0ڜ�
CT�Eʞ��ѳ�8>�m�g>,!
w�X�+�ĺ,�R(H�T���K��L\\Q���U��+߾}�%1�i0f���j)�O�b/��.^vX "z��z�G��ƛ�l����ut&,����FN���@�Y_ޏK��,��KnII�Gc,�J�'U]����x����<A�x��e�篫�\��-M`���e*��D"��F@g�tttLH������`G~�y�F��L�'���^s,�������"cZ�e�ju���U%]��{��`���������:���x�h=Jg���i<I$�r�mmmh�٪�O�4گ��� ��8)ѪhI��7��Ocמ��ר5�O��uY{I�d���Sީ:Fҋ}!�EEM@o�5�9�  Y�i���J>K���S Yy�i]}��03E���^!r09�}��*\-�y-��q##�.E�F�MI���J���~�F���L6��^�aܔS�-/c?�}+�����y~���2a�qE�;�#�FU�Ⱥ��^!���?�M��F��`x]*#��K�A+9R��B�U�ooeA��\<S@%i�����.>+��h��k��Dԧ՟S�QK?{T3��2�X;g�HN��\<��^W�JSV'T�_���p��,���摁�B�!�ȏ����5�.>���qlM����#��n�_*�xSQ��p���d��W��-7Y4���~�� <Qa� m9R�xi�ie5QB=����=�t��qEQ�
�<�B o7nn�i+=�p�ǣ��{��%`U��,��ɩ�������z����99��q�̼{�i`�&�x,��%Pa9 ������)p���u��n-��w�f��Wp��o/�}� �V�,��Q!�������-RWI����q߰��p�F�%�|i�-�9����8<��o�|[q��Ϣ���*Tߓc
�}�ػjN�P)���E1̔��F���]9�E&�����O�������sO;�8��V,.�Ɵt1l��3:�K3�R����ɖۡ�7W|DAa�OV�1u��x�E_�(���f����Z�^��,��8/~
�؊�X���9�Ġ����& $�F��vAF5<ϴ������_��'_5�WiF��>l�f�R�
t���I�V��F	/ԇ!PK���E�)���^�0�����a�xL׊�[�����t۪A��[�#!~�
k*��v�������g�
����������q<Y���-t�4y�cqU����QjT���F�<���d-Z�=�Vn<�x^.��<�۷�G7���(N�q������W`^������������*�Y����Mӎnvb��K�n��\��p]&'���}�<6�w��~��b6����[��С\�)�zQr=^��i���u�)����ٓ{/[���sF�	�4��q�D�a�g�����B��h�Bo�[�����tOQM�7x�k\��?ȷ�T�r�/S�Mci���D/��O��,���TF�O��%�E=ă�h�6L���d1Ԝ����_rl�?%�G�P1�����0���|Ի.!�/���T߽���NE��rnx�L�ѓwm�*�o���G>ky��)��GK��Ѿ+��|��|h����p�BLJ���e ���b�xH~ԗT4ި�����C�a�����щ7�MD\�����Ş�3���'m��%@�dw��
�~4?;rܮ�F�R�kʊ���4��O<]�Ϲ4e�47��k+��3�{◷T�I�%�]��N Z`�Ģ��;�\�ܝ�����_'勐b�f ��Ζ���B�P�������5*2nM����Z��Ջ'�-[d�5�q�w,�w9��]5�������-�O��IU�kuH3�C�����\$9�v��t�>��oJYHL�l�"b7�N6m��G"��>�[۱ިK�w���I�,2ol�E�#���.�L�,��Z�P��&�r~�^4����T꩹O�~9E�v����hQF4	㌛�d�^����������*��Խ<[sԈ�M��n�4)c�..��{�L���h��0q�����P\+���QDQ�&��x�5�.���Y-h�� ;�m}��f5hǄŰA���R�_FV6�F����-�@������|h+h�8\���=J�q���"[b��wu�>+(�y�`jS~7������2Ʈ�b}���@iT;��ڎI���@������8�@��!?��E�lc-�����v�+�� �G��u����3����*�rrh5��Q��b�G�{FK�F ��5�=�^.4�5��v���x��p�?��يHyݷ5
���!���-i��J�Y�ᮺ�	.�X����;m�<kv��:]���`X>�i~���Fo�%���9�7����{Im�f1����پџq{�6��|��tG��X���>���e�p�w�Wm��4+�QA��F<�I��黼�u�lY#|��2�\�s4�B����CR����8�󵊟D���'���@oprr��l�������Q�F�i��uB�\��w+�S�^7+�4+T�~�UT�n-����m���zd���	�MK��*����kI���_�9;ʫK��	N�?qZJ8s�S(,���'XK\�Er�7��4p���~�ν�0����Q=��C���p����O�B���������	��l�������$Һ?�κ߳�=�dX:X?��fo��Ϫp�M'����΅Rqm?���Tg�s̟��䚴�ғ'�����3��FE�fq#O�U9�ߓfii���2�m����ѿ��t�	���#����H��߹nOD3kZ��&�4x=�������7�m��:ar�O��	��Jzq�V��.�����+�V�T���*TO.Umu'��x�k�NDZ舠auP)VfV޴�����b�tW��Ek� �m�g.��ae���B�<���;���ThƸ�:�m��K��2��~[g.k^R� ����n�̅���i�{�[�b����5kSD&qU�X]���-�X~����QY�yk���v��X�ڔXM?jŤ+�(&��L|l���.�_:yF%���f/u��ed�����i[�7`�s�$�91��}�B����Y���bA��d�4��(Ң4?��UHd��q��!=�u[��9����.AZ�i�.�
:Z��H*"kwqA �$s������<�@��%�hϹ�Ȟǖ8X�р��������tSh}�X'�1���\LVz��q/f�*������f.��v��.6�o���(ۺ|�� *6�>wZ֦�D<<�������<����"������M����b_B�(�ͽy�#A@+�����6F@$߾)����1���!L$�(q$(d�"�PV�6��h�(o�(m5Dn��p+���񝳥��n;gf��ُ�V|�GgKGg�11YO��o�ao�Zd�!%�����0���U��������ޜ��wbI�yH\�������n��dVi��>�X螃�GMJC�G]��q���s.&����b~p���@s��@M]��z�GaV}d�Y�\x���$o#��r����".kw[+o��"wX:�pW�j�L�$� �sO}�y~��օ v�=<H�`�Z�����	�\���w�j=�;�0؍R�Q6��FA8zh�5�`HU�e�m��ܪ�L��aQ:Y���ҎKr�2��ۑ�T�d�8�L#��nA���Z=����݊h�������Pf|���N(M�i�F�Wi]�g}q��Ӥ�'rΫ���Ӣ����[���C�Q����(��Nu(�|�D�$��w���S��6"���{#�fa��G�9��E� �tv�:{�H&���'��G���Q3�։���H5���Ԩ;�!m3���k��}�j{cᄅY���?<=�WٷU���5$� �m�KJ`z�=`*̸)Y����Ma����?F���G��XT
"9p�C���$�]� ٰ�ϟpb�S��%
'��7��	�_}%��'l�^^Ssk������A�xu����^;��S��'p��z��z#�W�qB���
<)uR�tø�JQ4�cwa�ɖ8m::�]�r�H��f�F�H����;��D��^��)�t&��ݲk�z.8�%�]����ؼ��~���rK��B$m�	Nf��=�)�ō��ڢ�U�~���9��G�?�h�Qn7��+٘�!֩��!fS�@�<�>���>t�&`~o�34=m���4�V� V7���Ą%�E�ʫw���fc��f�T�0*e��P��5��[��8-��"}�]�B�rt����l6 ��5�gd	�G�q_p
����=��y����(�ء�J�5>�]n��g1pc����z�<Z��i߶�Yf�F��9�.��g�Mn+�HuP������Q��~��_3�;���@F7嘑B�3��Y+'YGfv��~]��n�W�{\.lsy�y���+޴��%��)M�F;Ĝj�r3�(w�<�1�^)��w��M���k�W��}F%my�fc.�7It%�����<��3{�zz�k��Kx�ޓ�C�A��V#,�)�	�Q��Y�;��A@���J�k����EM�ՎX�r�ϒwcԘ�-�Z�@�O�zN}}���
�Fy8�ܝp<)�qqz�W)�Rʄ'��941�����=L3�j�����(�0^rv����8��,����<�Nh��:�@�><2�%|4�t������z��m%Q�75q���k������%�K�(>�i�t��6�����Z�-�I6le($�RԸlT:5`��$�y14LW3����zŊ����Jzs�!�ڭ��i�k`�4 @C�ׄ�F�q-ɼ���T������L���B'���SY�%�m��yT	_'��6v@�~2��=�f��b�j�{�_K�v�D��<�:��y�$?�A��X�6P���;S�V*�mO��u%�9;�
��K$eM �'���\�Q�Rq���8����q�[��N�R��C�^���	�er�6����씌����^љ�
SM�!�p��$�����i��g����7���su5�Lh��`�ϋNsl�`ª��*|c�rfDApˤ:O����G����':;�ٙ��qw�"+B�Er�����l`1>�D&�G?��K��ύ"f��^T��7^̳�Ч�+cm�1�����@�>��?q�u�վvsӊT30����O��c�ׯ---����i �w|��P�bb��7BP˲�佩�.�&����0@F����<,*�\*��x(s`(,�+a��{A�i��0�?#c£��feC��t�%9��� ^�U�p�����N�F����K��]�G	�Ppߘz�Pu.�=ԧ��!L�AX=��6^�b<�o��6UC0Hݣ�]7��X�M]��t��QM���^�n����[�(��n�cY����.���?���׵�BB�%CGG����ոl�JC;�S�N�+�p�ɯ�����[_U�}=���ȃ�(-(�-�"�%����AH7��0�H�Ѓ"9
�C��Đ��{/�|>��{�Aa���9k���>�И#7>j��?��.�V��=���@g��U%,����
�s�o=�l��0ඞ~Y��>'U�褨��L�:&��A&��UC����AP�ZOk�����W���g< 9`�ed�(2�2�a�;|͹�3�2kR��P�S�:X�r��Dl%`�� v��`l�&�����%���J�����rUK�I؅��y8���$n�g��<�V7Z���sO�������b�`ss�>oRhh���Ժ�q\�:���J���n�Ql���K^1�؟�V=F�+�iVr#1���ʅ.|�g:Bŗݰ�\�I+6[S)���,Ze[�@�����L��2�q�2��N��RF�?h�]��!!%����N
C
��t����j���`��� �9|i�+%��:��<�~q���̜x���]uaf�4�}��~��^�R]�~{0�E]7U�[&�cW���
�=#{�� ���S�/Ow��'���M�#��E5r��%z�m�o�7|����{J^y�}j��2";<���g!�5Ri����B�]����5�~�}�w���`�S��j�$@��5d�N\�}���u2�!���r�c.�$�M�,*��=Kj��Y��N������8�C���S�C�$�_|���|[�;�u |�~\�y5"͛&E@.kD��� ���et�qԧ���8�<�*��4��.�9-��O_n�^����꼈�'sz�T�7���(�u@�n���G&C�����GT����4�gw�(|:(�h�E�D�Z��ݨ���'��,U�+b��˵�P7a�}^��Z�Vg3�f�,K�/��>:$��0]_A 봰���3�L���q��?&ߪvb�}�%iDdd��v��v20������%�G���ڧ�{��8�$�VM2�Տ*@�p����$�kFs�cE_pl��z��ʮ�Z/q��M����n�~Lkh�_���7#���6_�L3�3���_�9Û⺖�^g�y\<�1J�ȱ�͚R���ðE��5�3O�#��	�S8�;�ni,f:T���nj���F�տ���mY�n��0�}
�EdPp�H#P?U��X1+	��Nj�o����J��!l1��G�O�^�[w-q떦 �p���C���eB ��k2|����\'�`�b��Oma7?�IS1n?��z��Z;�L	�����W�:��Z!;������N܀���g�`�y'3@&�]�Ε�|�п� [l�X���I!޵ۢ8# �q#���yPD����PR�l��A�]�g ���CCZ��)���V��b�(�ɾQ;�z��Ip�N�J27	����P�� ��ܝ�\���[�C]�>��Đ��~Q�%OѲz#]O"��]#�O��4�Ҭ����8���Xvd��9|�raŜ<@7uT��� ��IQe �"@��^^�xߗ߷���Fl�[d��Ie��k;���}4\��/#��'XR)~ݎ#����� ��K�$���glq�����)s��O�&&&���K��	�G�R����u$}�>�����G�Ć�jg/��b�Y����tjO~4��L��2�S̘������A��c���_9칠W4w���V)N��G*��af��oyj�~���� >��lDo/y��)��dʵR\�=�RNt��S\7��4(Gyf0Q�s��g����n��ٚ�(�i:���v4�qN�0�4��|&6�@L�=ܿ��%r.p䤅@�6v�l\]5�̿�3 ��?�8�չ��;X���^dw�Q�)y�o���=HF�����#|�轸h�[4�fu,��;L��FdB�^��&<�e4(�n�E��T��EJ�3y�����# ���	��w�_3�9�so�DTFXd,�}���ƆNwe�x�%�t�O2�Q���ۮ+?
��M�aDf v;x5ZeE{���=w �xxx ��5g�lp���9�aT� ��M�RQI�Ƈ�r�}����7�u�R��&���C#��)�7A�9�k8� �a㠹޲��m��4I����Su+>a�+3�kʽlɤ����JTt�Nf�0f�-Y��u�bK�a-����UD��
�;��#�Zr�Up�wD��\�D�Y��	S&��,�(U%D����p@2!z���ľ�B�C��x�/]b�֙��j���(#�r;��W�Z��@���1)��<�`�/xGE�߈`O~N�K�Dc�t�h�x�E�J�s��R@���i��n}<�5ģ���"õD�����3�����P�- ��e>�]ls�	�.�+K�5����E~�;�OX����{�%3k4g��!p��Ps�)ǶZk=�����㗤�v$?�"�Q�V�؛rz:y�I���~|��2�W�1�@I����k�"韪P1U<"��>�}߀Td��!��PתN��W�K�F5�1׈*���Pϣ	���EΨ˴�g!�z;J�;�-k��r����dU�v:2U.�ƺ����q	�?D_N�����}A�{ඉɳ�������a��A�A���6����ڟ��7�:^?�lO�T�@�S3Pǚ�|?�^i����.H���z��d�����Tw��;Q�ŖVyt�ȸ�tP��Bz�d��Dl��)b`�iw;�{Q��G�f���UM��nXj]�b�З��dk�I��Y]���X�ks��O����pǖ���7�j�m99� /�ėS��---�� [f�bn;Z%||��Ѝ�x�çCO>U.t`=���<�F�|M��ښi�ҡ�.d���?�҆��r�=�2y�2�+��L:��������Z޺ő"��!�}M��a��\i߱��8n#q�><�����$mjMu��5��]�$�1���z�ćq�~���^Z̿4~7"�����jx/N|�O7ZK��[g�s��=WRx���q�ed�Qo��ۄ[�u���x	ֽ�0PY�ٷ.bT"u+G��`���D&���j�2l|�hT#��s$����l�&��n���T��\����&���K�<������{�������5�nV�17R��A�L�|<��B�y����(Z[\��R��QJB���TRf�6h#>M��mi
v�M2;褋�ܢ��``�A�� 4t�^׻��b�_�6j��q//�-A�M�M��^a�!֪e�3��hh�1���"9J�3��,��7G�R@Gbt,�p�?x�B"�v��Fs��b����G���'����{[�a5OM��1)D���C7KLHh���Sg�T����&�5u'���E���1�����5vI8ť`KK����% \��{#����x��C1�4�����x4z���zc[�J��~dmii�u��ש���*M�[��JѸ��Eqkj�P��Ƀ��x�&nX@2"��p��(._߷�Fjw�� �}�*�3�#�S����5�[��m��ʖ�t/#dc�9u¬7�&��oqKz�X��w�Bۂ��z��� �?�D�ή\ Q��[�9e�U;��η�u�4�T7�aM��9�rU��ر��5g%P�.R�'�|��^���ѡ2��w �^�C�e3*��j�˔�S���V�U����_.�U��sN�zԑ�z�V]�S��sLT4)|Qg<��B�^�l}��y}#ڛ��mGh1��2id���;u2Bϗ.o�Tm�Ib�JJ��ڕ|J�GT�{���z����������_J�#x>08D�����;�~�n�M�$���G�k�I]�S%r��fOn��z��=-��M�s}��娗�]��=Z��#�GmuU%���Q����&]��8��I�@T�;a�i<����K^z#?.�0�S]��/���}��y#���qv���ٝ
V���Vz��då��7@V� 4Fu��)vx/  �՚��������u�%p���V?��u����.���(&��Μ��"������<���ª=Аd�=��[i�j�#/��^��ʅ��;c�@�s���%���d@=��6���S�_��nY/K@/���l�N���s+�*Y*-�l=��H`0��;b_$Ѭ(??hb�Dg&�a��r�mx�PE�7��R�
�7r1>E���LS�q\����.[���5�ky�\��3�����S�X�.�i������V�}j�������'��}S�^��K� �#*d���,���+w��̼E :ⓒ�����k1�����i��'�!��J\�q���k�5�7��:>�\����Fb'v�Vq�p_��y��\c^����閯�K4t���"��V����]F^G>����Ѵ��\�jc�8����������@d�9��V\�~��K�Iۙ;:6���+�v�d��~f�n�P��>*��F�bg��m{��o���q�S�ҳg�9X�ӽ�/\*��g*fϥw<27�G�7���!-���j��M7�^g}*�wP/A�h!
��s-�c�slʕ���1�=`����L_�tp�p�
�_���1k�X����B��&�e��'H�[��y&G T�Ҧ_� �a�ت"A��g2�mX�&o�u�n�����
yq��V�!�x�Y]�'���վ0��a���Q�ҧm�]�	�[��2P��Z"S6t���<��(��@������k����)����͒fyYG�79�� :"���%(e���j��6W�V��A�"[d���?��oj�0�Km�]tlU$ѡ �N���(�bά�;2!l�Ud�l�(���֕ ua�| 5.�� ��s�X��`S*!����������}��H��0=�13��������C���^�0�C��v	�MrLj+��@���w݉���7b&sy�Nt���6I�x�v^DB�A��]��zn���L[�����с5��7��ߊfe8�Zl����g3��O(`�V�)�$(͙7&h�$��j�W��nha`��yO����t����S_�N|N������S��z\���������{���-F�y�b;�� �����P%�4 �[��A>��n1׊�x-�5�N�m��r����Je5ӹ�H�-��.r��Ƀ9�|-UzSe'�����Н�޾=��pP���<"�Xa ���f98|�2�(�`��}¥�ձb��ҍz
(��ru��$�Tu����L��"�Nxnܮ���H���	~o����q���I�u��D�F=�"���-�:�R)h����;zU�w,���l.>C�Wk����wu�@���`�'&V��$�'� �z�4����5;�E�"G7Cͼ	?�9(o8��k�T$�aTE�I���1��7ʫ�6�}4+Zn���9��1��`�;�i^)=�׈���E=~l�Z�@�^�߅4W�:d��G�}+ڬh-��N&� =�v��%s�.��Q��(�#�a�RՁ#>�b�f�s�z�FR���F�	��d��.�)hT�A:�(�bI���W��Ρ��{(**ඬ�/ "���PB���g�U6m�'�&�9pI���r�[�zJmq
�'G��B��̹�F��OrK�W����FB�\�sT�'\�q�-7��4�?��7����c��/�9�=�����h���^+�; �bCC��c{���B�VVW�W��^��V�i�P�5������Q!b��ˠ�ܠ��12x۵'���*ȏw�׭ݤ���Xm��\KO���x���p��B]ʊFG)8[�њ��WA�w｢'�!_�,ڥ�^�V|�v(���ϯ n����-��%�/tV�s�`:E�'��Nm��W^�b��ҥ�����h5����x��|.�j�{ls�V���!S���'Ԥ�ٳ���]����'W����\�.ߗ��4��kZ?C�<�}X���MT�F<k��Yt``��8P �MLL8��S�*j��4���SC�����˕kz#���p���E �0��FT���l�����+�Ic���?�*���a�E;=8J����gAH�҃���݊ļ�(�b��ɷ��n8����P��T��B���<<�b�~(%�%��3�^R��B���3|h������X*��o�׊ �pj%%}��n����0�'��{�k��=ș��D���Bod���Q��Z��L5W|��������P�j�6�CV��'7xF0�cG&�23f�<5�c\w'�@n�3-ND����s���8��F�X��!g��Q�ŵX5M��R|8�S&#k!_II�]����0#���#b�����Ĝ���q��cH�f_I�:2agP��#[��^�9�=2n>W��j�,L�D���稰���:��VC��+Z;�O�%(����ï���{� n}�N���·Cte}�F0Ӂɵ���E�=k@hٙ��������@�`�C����I~�%bZ	�De5�ӳp��j;1�#ur`��)E ���|fR�B�¢����"D7ٛv��G�����f
� ����e�շě�wҬʥ3�h���|�����^ʥ�8�A�Ѧ��K#��.�g��������Z��w�{�����:�l~3Dc���Ԫ�����?ٳRϗ|�0>�^�f�3�^%,�6{Eo%l���5�3������O�b�Xk;;�S=��s��s���zj�Z,��z�v�"r���G�����n�wq
�C<W�B���c��u��H%3i6bHmr-�3�m�j	X�?��4}kB�M��Հ����6�\c���G(�3�A�	����`ُ�0}B��ڌ�ho�^�z@�W�׵җhO��c��g0���>t�3����=�o��ɹ�fn�iTL��ߝ�N���Jn���@ �#p���<�h���Jm'�oǮ4:�X|S���C������iy�Ў�]]mP���!OMF�t��?s����+.=���uB%����:���, 1BY����q�c*=m�M����,G�j�[d���z>-�-��]�\]�3<���񛝀���rmWE_�Z?5Po���%ʷ9�j|6��|��"��ѽ]�z�^P�/����q�x�2kTB}��!��	�H�h�=�b<�Gc'�'2�z�~0�;�0����[���Mm+e�{�u�f�U.=��+;⻟�%2�	8��+++�{~v�2@�u��QO9eU�4e���-�==�6� bv���0�����V�٣2���1`���3i��#H�!���4�Z���6�(����)�֤߽�8���8A2~��~�j�o$<����81FJ:���^"���[kT�����,�����E$hr��A����% 5nL�*$���L�,!G�V��XD:��F썍��6��IW8�Ӣ�H�AB�]�- ��&�Rg��6�0��z�s�M�z����w*.�sk7WD*��t��Qd� }����ȗ��_��H��G�+���׈��@���0��޳�<������j.6]��M_gg��.�����|�ӵ~{��/�ܖ�"*ʌ�V��E!��m���-�7�O��w�&�4܆U�p�0Z��� <�ke�>�i	�,�[��gkF�qRd��]��چw����]�_
lq��90����J�=0^�����^@l�:B���_���a�ɞY�n�Z�"�Z��3��Cm��/����C��
[3��ː���MO��M{{U�O��|3}�t�n �8c�՛�eUo0eB�t��d�NK��A��]�֤�&�1g�x�>��Z@��"�`�hgUT�����Dúz���p`xi@["$(��6i�+)q-��3���;w� Ln���+/�Y��I���{��r��H��5��C<=�Yf&��Z�ͬ�%��{4Wp/��6ƽ�������$Da��a��IBc����5�h������^/O:%R����I`�j���֜��zz�5=9����[2��l��=̔�c���l����d�}�#.�x[`���>P�Ga�l_�#S ����9�
��G�{�*��`E���x�^լgO �	��������nb�Զ��Fм
�f���dԫ�	��Y��"��G�Ɋz���$�Dtj�w�uw�k%�� 3:d���Vy6]�f$�/���o�J$%� )S9��}1((��i�$��߯�t��=�2�XGG^ri;M߬O����[n��a�LTe||�`��zQ���(�S@)� �4��v��Z�u�����'�ydJ���4I��I���1�>{(T���H����q��x��Un_���Mne	�M�k@A��8E�/I�~x�C}>{�,�m��"�X���B<�29(�>@N~~<2y�o��^{e�(||`o_���K�ug?�oT����oHO�	� ��D���iNe�c�`��vuբN�����z��nKG��#M�Բ7"�|�.���t��]g��3؞5�
E��|!#	���ۼS����_s�@r/V&���ܰM����p�u���#+7�՞�(X�`[�㜉�	@�f��!v���q䌺������ވs�=�l�<��5}��Z���'^��6l@�ӏ�ٰk�HX��TT+�x&��Qw����RS���2w�b?�d*�.Հ�Cl��-Y2�{36(��Mzz�?5ï�u$O�[o#� ��� 7Y$z�:6��5P��i��5J
�>���%�
�9I�y�bk �}RNh�G��l4��:��R��e��C/���Pq_p�����i?�����Yu�
T)r9�zl���� נ��������biY�#�UX��R붇���A���D���3򦍒���@���I��X���-+Fߋ2m�/I�U�=��	� ����	���?�r"Nkg�0�Y���l�qR�<�{�%�&oU�f72���Δj�*��* �^8�+����}'e��R<ڮH�ۻ�c��Ѕ��l�ł���o�īh�Ǖ�h���Aq��_�4���r���X�;G�\�v�X+�n�}�$��84
vY��1&X{�t�@�R�!�����~QvK��-����h
�=���C���@K��FPJ�<���BZ׮��_��O��Yԓ�k��c����n֌:4=��hd�O���V<$�äTop{�G���]њ���rp	�������I1���VO���(��bˇ����9�N>�#�k,�w3�6�>&^��p��,�3X��@�;-.m�A��DȚ�$�V��.��PŲkW\��W~�A�庠r�*Q�u��f��Ml�ºE���IV�ʈ�̑Vj���0�3���!��l;S'�ZMS�R���j�OfhV'#���<��}�\�l��m���oC�l�����r�D����+��-%���u�o�~�ݨ���~�Km��ş���=+���>�S�7�b��7��������Nt�[�<�ǵ'�+��/<����P����A�2�X���ȹ����V���?��6��,2�U���r@{"�v��/f����#ã�Y vfZ0�#ER��f��`�qk�<���Kq�� �
^��mju�������׿W�VYw�\�e���Q"�o��E���N��4\�Wt���9e>��&�_�I�N��m��V�wz��7ʓ�w<�g��;q����,�IE84�=ux�I=�����Q���8��|Fl��@�Mg5RH(`�Qe|ʶ����1}�'������C�� sKq���)Ɛ�м9���Hبk�ޭ+���2��;��!�@�m���X�)7�X+��#ރ�T+��-���an}��z:�������ig4���VQC/૩
��+��/��Rq`�O�,k
��6��[�OYk�i�d�e#���ꞻ�͒���&�Z�"p-���!̫�l���&��ZM'� $d$���D�N����w�".8q�Q���
��R2�G�!<#�E�A'"+��ǐ��N�٨��%��L�L��f3A�_��NO��?50�/ӑʢ�lm;��LT��]�̷�5�v�Jس�N��Rc,>*B�=��|ʀ�R�/�-,��j�uZnZ_/�J��`_8l󏊻k�Cu�O��UOJ
��H��j��]�����e>k?
Kih��"Ǵ8���ɅV5�i����o��{��n�>��O*��HР R��BS0�������!���߳ ��)������c���C��-���}�鞵�ؐV
�1H?W�䁶L���i��g����0!���!#ǲ6]dJ���z�n�������٣�$O�Alc{��P���f��vG�����uš����d#�P�
5m�w��h���n�U]���a���k��~�3���Z�N�_���=bE�z����x�WO�8/�� ��l]t�@[ ���T��3Kٯ��.S��<e�������JD�x�������48�uO;��!�?K�{��wn~����PMٓ��*�\��Xx�vR$�kYw��x�J�w�&{w�Dw�(+O�A����>�m��;��q1�j�(��{��B�����(���u�b��Fkc��<�Vhj�P%�z�[/���A���ԋ��!�cLw?׉S,0�6o[8�����n͒<�� �~�.*�?`�q	 +(!�����������>ņ"sg�?e��N-�/��<��}�[^��F�P�3��Tz�T����٠���7"�w�N���ӻvǵ'�i#�GJ�H	���_̳����V;���R��^#��4�0��Y�H�b�vv9GohU�?�7Ɛ;��Ɗ�F��N5��ߨ�sP�/j� �ķa����N4W*��X8t�ޱ�x>�I���m-��	Q�J�={F��i? \��Hrb8p���e���P���`K�� k�[� � o ��[� �g��@aG�^�=OΗ6�&�9V�̼(��/Xb��_�D�:���ݳ��B�hu��{��~>ɷ��2�}e*l�W. h<��/@��4�Q���ރ�耂t�j*�n�L+����n�>y�\�W�j���Pzd�cnsC|�>���:���-���p��'҆`��鷏���_�C;Ya����O,���^ �Wff��Y\��D�PSYlHn��V�C"��A���ډg��:-���:���9�k�ٞ��oj*�k9�	D`K��N=����+�����x��x�:������4$.�iL��_��/&Y�U����S�����F�+������t��6����m)����1��>;�,0�UXRRK"���Y�3y��Φ*��È'�q?ל}�%a���,�}�=]-���YV��D�q�)/� �<
�|:&z ++�Vo��<ǣ�-�p~�����捍O����5�W��i��C͟�X��~��赔T�i�N���s��ϟ��b���䖿'b���'p�@A�.;���:���m,@AS6_�/XY^V�8������ox��o����*+G����Y�C����Fs4��߫�O���{|� ��"�zN8j�#�{�P�����j�}�F����	

�ON��F���,������e��͠<c�a�;+�!��_�� ��௷��L�������\��*+�Am)���{�/�'���If檪�����<�H�spp���w07����5���J4�k��F�YY�v��������������:��NVCqaaH�إ9j���(���Ç��]w0hOmy�����ݯ}����H�,//�.�GB|���e��!|���sT��Q 	�	�����L���3���N����   ����h�hKuh�!~@-�"��\ o	�엿�P�;6V��f@EG�FA(�m��es���('�XCK+$��,p�\�AAA�#kDw���^P��X�&gUK$�SQ\A�����ܯÅ���hmƲ�0��?��r�`[W�8gp��37���C7跞)p�����U�����>���γ\{�H޸[Q��v'��oj����o=��wS��&�������=�n-ߔr���"K�~�bٟO�L����;�s�����W+�@X<�i#��9�P?1�N�cP8�*���6��n�� ��/�q[�l�b�_�]�����<�����54���~����,nթV��X�s[Z�V�+aj��T�<W�S��hv�%���Y.�'P��������L{�m��8ׄ��yDm�/9�\��R6a�E­ixh"��5}k�̰sWcB����f���ס	[�t�Ԥ�%7$�4���4E~���9\�"-L�K�h5u �j��9`�F7&��3|���0��v�ױ��Nv��cw-�����q�I��~Rҕ��I�Q8��v{��_^	��x�BR��{��L�$����8+�����0�u��e%��`�Rp����zn�n�@E��eG)1m�������i\�#��(��6��@q�ݥ��;��R�O�Ȩ�l4E	�ye�]4��1V��Ox��E���m��2y�(	S��FS�� ��-v���,�z�ܠ�H��_$��)� p˅�o�����w����	������b��)"	��E��F).!b�y�]��O�u�=�#>G�);�S��5��:�I��c7d��m���_��η4&{h0���w#B��:l����K��<<<��� }�4srr�z\
�ܘ�:8Jp�LBId-l߭�o��>4��\?��K�$y�����8���P����j��t2~�NG>�Q�"��<�����Ԫ����G>�g ����LjFݳ�f�xC
g:Q���1{@�)Y� ��6��,����Ҭ�x	�h�C?lg�7j
�TNE��8M�9���ic>Z%iT�D}O��J	�9��ތ�]����t%�۷^��K@kxt%�>�
^*���2:
��� �PmD
����|^��b'���se�eR���'�Q������0��Y7��]<He�ڶ��%K�L�T��۟9��ok?	.(ѯ��_x_9���h�a~��-/�V�mޱf`���9���Ƥ�xp��@#-���k���4�Ż�ѿSU��!���R�נQ&լ��\�Y���[���b���{���������+/K˧�ۋ�@� ~�{���3� U.ܭ7�qY��e�M��}���#�����Pb���/��պ��5�4=3<�1�^��E�ZyTKD��Y��k�~E���8Vk�\�dg������
�;GR�"�:���`Q�{��*�v+�w�L�N�����DWJ�4iۭ��j�J�)�1��0�j᧥����~z+��N���KD&rЃs/������R�j1�N�{s��K)>8�Z�g�������q�J'�W!�KB����/��UXN>V<����ɸq��P;�:%I9%�i�˪̓0�����r�G�F���7{5Ggt��n��jH�|{�}O������ ��g7k���4TUo&��^p���U���w�����D������3f�S�)���/�������k�B�;����f�<�=����0�y�3���w*�{�vZ%��������>�\��V?+{��5��򇲘��jhzl-�������2�d{�s����y�uޣ��|���'��q���,Ͱ�f��j-�Ct+�RˢU�����a�Oz�$<���R�ec�9x��0偬c S��e��{_�R�?Yb����I��3�I<=Z�n`Ps*����] #���(��u>��E��zS�{��k�����NSLq�텛�_=��zs����w{��-!!q�8����dk��'��|ƶ�f�e]�b+���)�H���:���է�S=""wF�����[߶��?T��j�4�Y��u%f�o�K�^������<��t��q��[���!S�E�J�\�Ͽ�����/�����n���#�R�ae��fV�BEK+H��ԝ����������0;���['���^%B�ʌ�G���>�j�ϊȬL�ACW����n�wE]��t�nѲq�y���/ɕ�"���wŗkh��EЉ|N	�egUp����@�>�ק�>�����w�Q�8��.wETݵ�]-p(3ߎ�t�?�x����%1�ؽ��;,Ȧ�x��f���u���}+���t�9���o�]�JW����ۙY���tt.(��JQ	a"��Gl�%�a��Y�������+ (�Ɗ��T�]��R�C?�9���|�]�Ue���nz����k�Z�9�S"8`�-�8�%�Y�z�����y�B|f{�M����[�M�{Y�y��9��W�e����h�sAfJ��U�Ϻj���D2�}�޽�A&h_�	
���޽{���VQ'��ic�F���_f�э����O��e;��^��#�Qq�9�)*�V�����C��,�����c3^P�/�
׸跻��dO�Д�u���/ɤ�ۚc�=�6U���5ut����U�H̕D!�ּ5b3ۥf��4i���y��k�ќǜK4�7�`�E����P��mP��fpT%�������	qu#[d^������ <�� ���c���!�xz�������:}���~�ue�y�B�c�h�o��
�g�������r:x���ZvN�7�s�E�()�
���b�����s	������[a�"$O�kT,y���{d1W)�)�Ho�d5ɉ�5���8�ZtZ��mf��[|�w�Ia`�"��;ˮ��'R�m����'�7'������6/�����-�e>���O������P�- 
�jrʿ��^K*:A[cQJʼ��D��2.�JU6�M]QJ5eQ�#-Q�e�Dԉ�e�.o5���;r5�!������W�o.���5\���7���y��$��^dq����ʿ/����*$�ɕ4��ҷ`uu�)��m� ��'���+@���.�+d���DO �	]Ee�*�Yi��G�������i!��r��ȝ]O�Ŝ�����Uei�a�a_��D���d��4d�^a?A�#h�b�$$�]XR"}�i��r��ůA�2S�[oO�������Cg��qF�b��
{��m��:2Sζ�ʻW�V|7���{T���ߺ9S]�#L!�9��-^�*S{�>��j�#����0B���Ĵ�=RW�z�����O������dɾ�������O���,'�f`�g��m�U����{i�����\�x����EB�)���9�Ⱥڋ0�w֯���3�Ĳ\�c�f]f���	�OGy�<���Gh�<R�|��_�ȋ��,���47�ĳ D�@�m�{�}����-�C��ؔeZ��a�'6���ڒ����|Y�x��
Ӭ�| g�"s��j�8�������8O�L��ޕ�������i���iH��8�o��E:��W�#�Yd��&��=ʵ�{�15�I������������ª�5��SM����ݻL�-E�� -�{(y5s��%��zC��y��3����b�Ɠ�V�ד/�k���M�Dڴ�i�ǚ!u�WDu��u	�察
��i�t�����ۻJ��(.��=��
��o�H�(R!7KlR��4�p��t{�ɞ���[ݍ�<�Pվ_��em�f����6"�XD~>��k�9@��prp<24d<"|%�BIy�K��
g�I��~B��`��\���~�eE�U<Պ6����3ۯ�c�'t,V�o˒�|��B�~�v/f@��^�1t�rD�����\ĸIx3Q�����e��?~J�'è.ob�r���kʗ�\��Mk�x�b�@��}�G?L���11ީ�z.��MK��S�`���7��k��K?Wz,-�lnA\;Q�:��O�ͺ������IaJ�;!B��׏~=�m��9�r�p!%(��Af�G�Ї�&�W�'���K>�+ڟ�zPJ&��x��溛�#�Ȳh[E�[]��[�7�i�TxIik���[Vk��$�e�A���Q����̣�o�-]�=蚎f�/�W��~��={4�y0by��(5�ğ{?����}�I(��}�_KfY��0����5�
B^ ��c~>IJ���CH����NM���MY7�yۉx�cj��̄A}�Q�_������!�xJk;�u���%I�R���lH#���D�Y�K]8��f��C�|�9��W��e�v�6����9`L�X��L��h������b �]�	R}��o�6z����U��R���Ϻ���yz�"pv	�H�ߠ�485�ٯ��敤��8xxd��%�^�
��#'�[a/��Ǵj&}y�lS;��L.b��0���sJ�l��FImMO���vI�>0�:G _��-%}�G����'mY)G�9.��;��hM�Ic%��&
T�P��m<5��V�D��d�M�+�
��~"�c����{|�w��,-�Î��[]o)Z����)ۇ�$�<��C{���y�,n�� �R���-��*P��/��ԥl�}���^��տ뤪w�����y�m���W� ��v���j�V�����{!�jg��p�2EE�o%zu�2�
�ߖ��й�"�5���3���ƜI��Y��
j��ݷ�|�N�o�U� ��1�p_;] �������L3��S�Y�)){�m�U�B���1���ju���V�)���?;8���~Z�٠���\@ ��d�����܏��.`�ZV��x���\��_:��k�����jh
�����CoH�Ժ����uh(Y'�pc�顡L/!J�)���5v�����cY"�[�4IS��%�^)��6��3PL��ͼ+ۢ��xP��?��׵���z�1�C0wA��lf":����Đ`��9�QW����S�R��e��9��ش�"�L]P��4�-u��\w�#� L�2��T��$�k}��X���i�Q��9�x�����/�g�-/��wtv>�b�I�#�FcD��B���דfwf��vQa�NS���"������c�=��-�f�
��bX��� 5XP3�	S������w�Λt1U��M6{��NtHH���d�z��8(N]����/p��Z-�.?̇\kT��2,s%#0�i���z���l����N��u�+W(]�ZV羸U'���1S�w��R����xa��]�ОX9b�(L	xz�3-�Z�:���=��u��3v�E�P�^i�|t˥g��>��K_�8>����#����=]|���\��36#������9�����;N�O��X'��,���c��&Ů�	#_�(��;~�A���p�Ж5}���~��1	t<����2!���V��%X%Z�bm�GlIn���b�����ȳ�?N�X�-��k��Sqñ�ۤ����*��:٤�b�Μ%��g�!���B��9o��Q��lR�I����v&����#�0�������΢ϋT��(
����]�'���W�c��� #s3���gq�7�uq�(����wUM�=��'�E��`)���������긨���A�CJ�F%��TJ��;��2�P:F��C���;������?8�}�^뉵�>���\r�z9�g���f���0������,�KU1M�X{^|�k\������~�AL;dTHgb�����/�-1�N+�~�D���R�F��xK�};��ײ�ʰ-3$<��NL�rz~~U4��_3�Kwމ��}~RC���7�w� ��?����k|,�E���	TR��pf��r �K�}EF��wQ-*���F)��lug��K�܍�Yat�
�8�LL��]>�� ���G,�x���߂�Z@�<�4�9��W���]����8�Q��0��I�����U�h�z�؉7`����\=N����M�5Ȳ�]rh��d���PYT]8q qp�:u"���>��N���}3b�|�S����u'giG�&I��Z��}ȵ\��b������C�:���r�����6s�؁'Y�bA�i �6	�Z��W��<���fo.;L89�ޗg�?�yS�b"O�0����'^[WWn�E���j�EB�F�����	~rjhxE �s*rb��2�$k|.��{����b@ԙ�r���ҧ}��`�i��xG�&��#_Q�x������|�B<��Lg՟�Z�����	��8����(����M�)��!�Q��ch�z��:7M�ýp3j<���x��T�����W���+7���j"��f�W��m�W�\7��m7t�����w��Q�k�$�v�7��xY�HA�tW�˨Ev��HCu�[!���#���!��~�+��eE���W�=�j���Q՘+<�9v��9�� $?�N�v)����$���A�����ŷ�&�jq���N�s�^���t�Ղ�z`u�Rp��?�=��S��qU!��{Sj��e�V�k�A�j����#{`��_7�r�هA��ά�l�x&R�7 Х��U���H�pOC����X��t�E��ן_�����F�Z���/���yыɟ�3E�=�����g��������D���rȍ�N�p�}+�3�@�qNif�Ә��k����*��v�"�#�d�!À�+k��@9%��¢����G��� �nǎ��K�%]OҒhܰ]v�ClLI��9�UǪNPd*�!�	f`xo����)��j�ow)�}�0Z������������`�G�DZ_|&���69�`ܖ�c���oԏ����׮� x�ʤ`�����@A��ϱ54�����R��%G#��­�S�FE�A�����'J���b-�a8ڸ����Y@Ff�)ī�{4�.y��|��"iŹR�c��Jm覈�N���ؒ��s W����I9NH�e���=��SW�r`s��?�$�'�Irer.�,��_����IiiQ���ii�i?�p�l�������X���W��!X%o��D��["e2�	e*$��K���w��G��I��e�t��z	BV� -�j[��#*�$��uZ_����0���ݕ�gë5R8�(�UL��j�(�?�I�9�Su?uf_�@6(LT}�����E��op��b�e`���2��q�E�ޱE<@M�5����� �k�|?@��8���<J��ȁI"���D6g`����\&}�W^1���X�&�Wy?��j��I�z��H�����9�T|�y�y<�wVd����Mp�dT��=�!f߬똨
j׈����]������[n�G9�ͣJm�lr@��A)a0�e�Nu��H@���LV����/F)N
�
����բ�8��׾:$��!E,�����Jז�ƺIݯH�����閄�I}�⦷ �t%]���n�dj�%�&���=!�n^9Zʉ���P&��g}�|-K�[�@��+��I�=?l�V�1(g����c`/1�L��󽘰�w�"��WM��1���[DkJ%�$��g
a/P�6�do����b�u�>5�a��*����~T��a�ogs�y�ʖӤ\�@JN�t㐂v�+��ʤ�h���A`�[4�9�M���đY��]�!)����P֠��aϱ�T�4��G��U "���~z�_�`j��@m=����]z��c��;��ǂ�n������)���hh�72��Ѕ< Eы�	�4�{	i��x��$��+����V��*r��K߾�-�'#9�Ÿ�?	������H4����DQ�5���mf5�~�tݶ'n�XiF��N�6�����lR�)I[Z��]���������!*���~W@i�@ �]Pڇ)�'I-�1:Óh��WEK�.i�WZI�>#?�!�"7#x�
l5U?�J�i빬j��2X�{ȟ	���i�N��>���T�a�@
��֓��1��C�T�ꈦ��nZ�y��p�Wt�����C�:�YYh��x���X��$h�d&{�Nqw
�RtZn�|��Mv�UvC�n�"��H�'y��������@S�uJ&�N�[-t_�x"���"S�.U(�݂?-���W)�mn�����������k��s��N������44�`��Gb�L
(M���I�u�'����7�����cn��fD�zVM�"1q�[d��9*�o�dA}T����B������p�nu
�d�*λ�ºո�M��1X�����!��A?���W�kb�&�``Jɝ�M�ZO2Y��'����[j��]���>]�m?Lz.��&N�*j����Un?+�]�Y�BD��?���O��X�u����2�ֵ3ړ����}��ʔ<�����`P��q�q?M���)"�G>���9�}��$L����(��Rz������7?Yp��cp��C��`�J�`'*K��&|���|9�Wd���ٽ��{���]�C܊�Q(�e�ζ'�M~0������:ܐ7��IL^^�\S�����8�Z�Q��F}����i)�p��qkLfe{�g!��sf�tA�D#�g�z<��#���b�u�6�4��%%����� '�c�ꍠa�}�@{��^�D1G,��H0��a(	�Ltr!�s�z��*��"$�c8��I�'&<�H���iC�iC�������f��g��j��\l-��YiC_l�=P�FSt�P��f���	��f�!�\o�����ˑ�p���B�w����bl&��VT���\6�\�����_3O6(ZM���K~��+-�P�C��g�|itK���^��z���Mw0ڼ4��O]�O����Ǔ��� |�Њ��E�I+���9�����eZ�W�­���V��琏�T3tќP2�Z�;o?�����5�D|��̀��#��Z�\�pp�0�"`�H@����RP�������W�����e �jz�$��!Dt��X��e������������>��:n. =Yax��� �����n~�P7=,����p̄oU����� �?�#v�?����x�S�K��ǌ�O���{�P���W��|哺&VO��:{"�s5i_��^8����s}�H)i�p��1��Ƅ���n�1��^��������ff�O��%�� Ҙ_��)���V���Mzv.�Yh��,���}j	
�Nͼ$��)��^�qM�Ɯq��<��-���*>HbV
�^A���잻�D�b)�I�8�! i�X������s�,��h��}ʸ:��`�b��W�n��>`�λ�x�8F}0ܫ��Gy[Y��Fs9y�-6�d��@��t7I"lDB�0k�
���E�Y��;[�&�3�m���/�0������=LǱ󢹚S
O��C�'UE<َe>��F���UVr� !��t��wT�l�-�X�1��sd��Ao�MG�X!��r;��le�&�3]����-��&:9c�jD���Yfi�U��B�r�%����o��K���^Hym/࿖��� 5yZ����L<�Mt�h:f�xh�U����>�ӣ��]���Gz2����8���;T:�j>����Z��ޫ���

n8�gffTc�g�M r�9`j�/5�*�;g��,�^������%�n��#ב���Yg�4�f�]���\@��}������w����F��9d��ĉ
q�����B��ɤ6/2O�@:�U?���I�4in}��0P^�S�����/��/��G��Y��+��~��ZΥN�A�X�Q�˦��]*@�s�o-��וNYqd�sAE~Rh6��i͚�HO6z=K��p�d����v�(�US���2qܷ����Mw�a��O��g��j �/p�4H�7��d�Q���r�l��Zo�_�'��v3� ��m�@�4x�"b����j��<6qr"r��~�U��PGZ8[�N��4a��P �� �Y�#�� �n�֮��Zg�����|>�~��q�7z2�d(��EĆ�+c�{�ړ5=�'�Q�9�3I�w����-Tb�=!�x��ĸ����s��w��-hmܤԇO�~a�Ff�&6-�D�(��"�t�m�wc/�2jj���^6���y�G�dq�po�+
 j~�q��T6F�=�(āÞ�!�g8�O6����I��c��_�0�L�Lz�X�˲J�[�e���2\M���aք����Өyt6�6�Ǥ�[i��c8�j�(0��x�@~6�M�2�}Q����hJ�ƺA�xĊU����@l�θ1���g_sG�UMaPq��s��v�S��G� +�]�/o�6w-��/�l�|߲?CJ�4�}w*����n�C=Oy����eZ]_0呐�;c�Vz!d	B��Xfn���3RyY� ؗ��a�/��{֜�fu�%�F,���Ђl�I���;3��	��~��������М$0���W�Y@�sB���rcst)}X���W0�����s,ʯ�䤄��# 8�
�����췳�J^�7�2X���!V��Y�mͶ�v���X;: Y�����a�떵P>����<{{��e:"ޯ�'~�
�	I��K����zڳ+T[<]y��r�G�5���D^:F�t�40	�0k���'WK.���)��;L_�J��=K`Qz �J��ڃ��
����xA5��r�Skv1�����bԇ?�v��IW̄�*eq�����tw�b}Y��S�o �_���]?��}g���@H����{��A`B�	�}�S���L�K���
�"�����{�����R=Yr����ԡWoP)�Q����/�Z��.�ݲx���HB�%
�@��؍%E��ӄͷ�.Jc �����X�|�vy���w�r�a��c8����y�&~/��l�7u'�S]*�%_���MrK���p�r�zLe&z�Dׯ'���Y��=.))���j錦6��A�� $	8��;�!`����=��v�`}j��J�|��q_Dla�r����s��P�Px�ڸ��#�s�e�:�{%#�	y
�mnd��GYD�Dhm_{ٞ�9���<0k�J��M�)j�M��`�\�����e��HA}�'
��ĺ�2xhN4W=���C�H��@�����Ty?,o=-�h�����+�vY�����-�8���ҊT
���Y��G�����Dj�/����?��őI\�g����?���&���ؗ���X�/�vP��u2����*�;&�xx#�� ��c�S,i�R���-�o^�n[CY% U�S����WYm�=o5��
���-�Ơ�B���3<ե��ԝr�Hf���������*n��M�1nv�*c�K_ˌ`�~jީ�#Eޡ�4�ƽy�����t�C̥�c���5�L��z�C�;l�7v)�n��&�վ�_�w� ��(O�0P��P�h@�0B�o#��*9-8��1�F��
��l�ʘ�5m��un��Fϯ� �,��K� ~l�C��[�?[VxL��n��q/,����x���~���!��4����aW�:�Ô�v�����X�� `a���-*��Uo�? 4H��Tr~m�h��v&>ea�b�-��3�fF�F����Z�XV�2O�F�Q����,<> L��	�o@�&�'/��6��S��a��Ao�>��6O���oH��І�W��o:β�x:>��Q�>�
d�4�d�!$6'����䏌�G+��K�h�?\}Ǘ�i���PU�H.۵�����>;/z,�|�	�V#
��=��M��a(B�q?u��((��Z>ʫ����/�3?%��,+{�T��9�1�q�.@��{aa�����@�2�"��uCY_Ai@j�������=��z�!<��4l#/T$��}�^�k�ͣ:W.ÇJjo?G��b�=Z�>���/=nWv>(�p�e��R"�#��O��\i�E��*d���5M�q~��0�����o��̪}O����MTQ�w�t�L2ϛ���Ƴ�]DٲR��H*u�U���D�Kl��P'���+���鎔L�N2 ��Q�_���I��%~�=��L3���--4��9���GAA0�?O ����t5�k;��G�qTK��^�k����b>Sܥ� ���2s�e_��Gw[qrr��oO9��I|6���P#��B��!���{cc��h��"��o�^L�!�1�x�6��P�r-�nʭ��/�^Rs��`0��.=8@빴((�~\��IVE�\�ͳ�/���eƸ�^<�n*3��ڏ/
޹64H���d#�"Sw���w��p}`=�^v4c��/lohWRP2E��W`�T^�c��D�?�`�.���]�=�g��48f�����S༂td*�|;�!�s�ykp���M���=�[��"F)�l����"��8�@��*�i�u67��5�t�.�}���8$DK���#kv1�	b����GKB��~�mg���&��A��csF~*	@,cOj���L �?��Tʡa�+Vz(h���o����r���Aj�����>��M����R�_��^E͑[Jy!N	*;Jd���	�`+� ������3�_�w��ޑ��eH���hc�� 	���Gi9�&b���WN/�j}��Z�����SJJd��u��#��ih�/
�5���o�\s�)��]��7O�Qx�l�>��{�>y��hn�@��؂��?����w!N�~+��F	0��d��<Q~x��n/�  �Il��
'�6,t#���O��HQiF��yA���p����T��SC�����P1�M3��cG���V2�q����/�w�FffzQ�:��ӭ1�x���[IJL���H��A�ݠ�̴�Pt��x)�x�9���E;�_�����#ޑ�^�; �$�!� ]�f�1����{nM�♊�#pQ�P�Z�3�o�Ҕɘu'�a��[�X�B�qǟ���v�~��B�T#��E=E�i�:��� �/`�|_�#���6�>�����(1_c�F 6���2c��vؼ`nnO�p��&��r��\X!`�޾���C�hϠ� �\���l�^�GIt�|.66p�;�x+鳕�:V��ĕj�	�b���9o����ﰠ��޸
0/�k���U�0Y%粦m��dT��Q���N>��;�J�ME�+�}���ո�S�/ՂJI�h{�������t�����J�x��G؆On�����ҟ��\Y�}���/��NvZY���cTv!GrJ���|tY�5.E$F|��)q��{���o�p$�C��	��Ce��̻W�;t)���D��1��ґ:>߄W̖����٭��I^��U���!�_����D�d��.�]U��Za�5� ���H�l4Тk� ��/���4N�tA����U^G�h���D�_�T��,��(��;�3��O�1�"Re��H�nn�����a��:�TY������=�_��z0��YT~C��<�8~OFN�w?�s�� ��}.�b_��]�hǃ����5��ZD<��!�l���WUx+�t�Hp��D�̌[�#<��L�5�����>X��WJ.d<�[� ?���TÆ4Ṃ3f��^؅}�B��F�t�[o�ܾ��:aQ�)>Ⱦ̜�Nyſ/4�A��q4g��,f�P�ł�# IL˿�.�<33��w�hKۅ�/�(HJ�l���$��͇�8o/:���S4�`'*}�sWlY�!!�����o*�z΄IO
��-L�U���kBQ���Rۦ�� %U\��U�������J����q�_�����A��0��"���tdc_�=	5l�	<��Pa�h���Ât�b8��>�/�2z���9XM����e����Q���v��M���L.d�@=����4`�⮮}iG/E�5����-S�/�� ��h��W�v���H�\ �)a_�9�7<W4
83���;:�]���P޿A� f��ޙ���`N�瀩�lo� �����[�lPb��$���-�����!qbbZ$�ߔ �{�v�,I��#& ��#e��d .��]m���FȄ����z������/1�G
@d4��3 �(�D5}wq�SE����PJ`DG}� ܼAl�`G��/����!Nv��pynv~��ذ�}���gn�Sl2?-oO�YAgO��PP��c�z1��Y���N��A�~˯C_���&�?=1rh?��"�H����]���v�FOM�L�\���_�~5o��E��=����̢�!��My4 P��ֱ�$��3݈�B��"��O6�<jڧ;0ѣLv���9�qC����+ki��I,U�~�ϡ�6U�ܗ5����Exݵ���V��]?U0J@5��d��;J=��:���k/��M�<`?*Cd�,�k�$0z>�b�D��]*k⽃�" d8)�!���!�C5X��<'V�����n�,��f�BQ���0�~�����H���=uAzJвnXzŴ|�c��p*�)>�_��.׾�Che�r�v���Tl�kx�<� ��f�s/�Ũ�3C�ݾ��ւE�+gt8{A�R�h�*It(i���$�1}��xm@ʇ����V,����>�.@eL"O\���F�s�8!>��ϜzDѲG�Ee �T�S�������^���wo�d���=?DF�})i=����J�y��N{�������u�_������V؝#�iC*���B���Kvq������.lǨ/x�_7@Vg�j��tP��s��p�/_����M��О�܍G�K���1��ė
��5�� �J�'Z���?ܽ�4�׽G�lx���A%)ˏ��U��H�9���W�G�.rh���9��>�9�� 8�ǡ���b�Ε�D���c[
Hvܛ�.��%�U�����{<^:o0�����y1�����W��	�>����ͼ���6�-l��5����;6��6�U�D@7r�X4�ڪi��M�
CV ����?s�ܖZ�qFܻ���d���`#�(��Ξ^Y �~�#�@�q�#��X*R�AǞ1�D�^Ķα�eP���@�cf&�Q�D���.V��`�;�E������'~�b��ܗm�����'�o�^��I��yx�*���Ȕ���=�ѳ�}����Q'����j۳gP&��\�,?TC���V�RL���+@�d���-�\�_u��T���*S�w�6�it���Y�~d�^�?g�5����}��o�ɼ�p^�rm������;P�f| ��0���i�D���qr�m|���?�1�;	ĻRMÙ��3���XU�s���J�������Q�ß���ˡΨ�1��H�����1�5��a�jN��F)���7�,5GJD�k�d����
  �a�t��V��.��CS�zrb��X�~d[�3
 .��<T�(

#J�jL���ۨ�ԕ�04��G��w� سl�qzIS�w�٠�r�S���	��M�
}������R�{3�hf��[:���������h�^��������0B��̒7]�}Z�bM-�K���l�9�#��G�O�%�Mm��]�_$n��1��.���:f����:kj>���{U��\�vmg�I�U�ؑZ���ğ�<�6 ��k���DOk�#(�;F�] 	�:����Z�9kK(��c3-��|@��5=��i�Wm]� p�V:�?�?�����f�G~>6�E��]e6����B\�)���b��\�Q��k���t��X�k��'�	��� n��&�&~2u(O�+9���&�qQ�����g�kJ~|�s
��2�VLf�ש�֒�ƥ�����Y�?S��B��G���F-#��X;��~7O�T�7�d)�����[���o��C���
!ɱXv�љ�!I�J�a�񵄀�L�Э�;&�	�"Jw�g\���b������I�ܴ���vX��Kg�&U�̇,�{Q�lN�Ԍ�X��{�=�kx8O4�d�/$%Z}���4�a+���]���|@:D��<� e������z���:�2�=!��S�co��|&SO�+�
����XUmrhSu�����.A�6FDhA�A���"e1�OgwZ_"
�3p�\d��|�_�/�8*��_���J݋�2K�%{a���8��v�u�[��`&�/E����\���;u`�e�r(�\�-�(����op�l�{x˪���O��q�,�����x�*[���_��������C�:��()P�^����~�h �>	
��C*�)k,��Z8�l+C����ijIk���k�=@��K�ay�C =P�=nX��2vc����,��@X&u^j�r����"���G�x=���>F�,s�&�����RAC��U�Y����B�%�{��P�D�q#X��g��SN=����u��8q������������y�\Ũ�W�e��U��'��o	@�ii�:���xD:k��[	�<�#��}h�Wx+�-�=?�v�L����(���3�� �hI`��D���?s�F�u������k���{ܔRa���$,�t�}�K�k���ʱ�$A@�V��D��� ����q�.�|jJs-}�����M�K狡���2uO�ߓl�FT) �Qr�6�\��v��� f�C���!���˩%�0��`rKd�I�;���e�����)�,�u#k�q6���w.ϸ(�dp�wR<�v�s� X"���#��Г��� �4�HR?$�[HH
ֲ�*��o.,*I�eV6KO��t��.���ELdU{@�2�i�.$�ԝ��B���t�����=��˨}Vz&u�1�J�Kª~��w8<�E� ���w����E5
1-��E,�bt�OY���۴�lAV`L1�G��X�֏{c��P}�5�hՊXOZ_s��Kql��
�5`s4�9��&���_�j����)��ȃ:�Y�꽪��R� G��G���L��'���Ş]��=N�:�}~�%g��%9=҅�96.s.�E��8��i�E�[�Z����?���7�5���g	c كȡ� ��䀿;�%�S��gR��y;��!��WOY��:�7����\o+NY�����LU���ݫ�_�&���[���c���������N6��TY`�3����
HL8���P��{t,�-��w�-�/����~~N�YO�T�j},eϹ�s��,̋�]�}��7���;���]���P�m�s'H�{#�����1�?bEz�xCrp�ܰ�d=~D�qc�UW��=*�*�s5��/T����m\�x?C��/�a�f���d;��N �x����.	u�n &�DIm�wCɪ�F߸("M�r����~��!�����:��
G-D1�I�r�4�xJ�OH�2�Q�b��ț��[��=q�
$@��^�' av�o��L�+Lw��=��;ob�	#e*"7�����P���]-�*����?�(��2�ÛH��B��X-]}��&dt��$� ���a9$�w����Q���-��`�����H4��~��X;�fߕ���Ͷ�"^kR���m��o'U�%��W�Y�RЛ9�}�:�3ts���mbI��J��N��,���⇉]*>�q_��x�G�3�����̻=�<�f�gÉ�G3����_ �'�E|�ך̜oL�� Xĭ�zE3[.���E0��F��S�ʉ_�	PCX�*�D�\������y�6����)�c�2xKK�ZW�����?��D�����g�g"��G�o�,6��d����.(���:�Dv���z����Q�1n�N��|�¥�p ƌ��]�ݫ��h-�z���wɳm��>[W�w����,��#~=��p�L�sO���9��&Ou-�v�"�_m����MO�+Bz:-�P� 3}Y�t���Fy֝3Ӂd��
s<&���䐲��p�%���=�W��m�1c��LQ�R3�I ��F�\��G�@þS_#Q��Tx ��_DY��`�ϣ�ܯ3�\K����rp��w��ڡ�A��f�B��"��C��NI�����'U�ETӘ�Bȱe-?��Xe\�h����_	�Ӂ��\B�7���a'���T�JFT_�^\��T�/�LK�yJ��k+d����׿�b��w�/�y��Hۦ�-�zh;��%���˽I�0a�β�Zbn����h���O0v��PO�Ǵ�(d���,� �#�,�=&�օgZnUZ7�&#O%0��vHd%|��y�"mC|h<���������l��L��y�-���\���aIr~���$ �6��<���}�f��=���g�Ge&�?&:��:�2Gd�$ �O����.�]��3��U���#ZǢ��K��/N��u�������Yȭز�7���Xb{B��^ƣL9��Y����S��$Pi���ا��� P������{-*����Y�>��6���A�P�x��b�5�u��Z�%A-Kۉ�hSb���&7d�s�.Cz��&E�3s��c{FU�Љ��ӜR����ʅ�嘮^��)��=�C�7���M�p��!��@�B�3�e�S$��������j�z~�뒋&���w�Og��rLty���@�/������0�|��]�d�F_"�@ Քή.~~�##j�w�c��U����W;.����g��t�#I�����H����]a���m���5ɷ�j]�%���r���Xي�aݱ릚*K�y��4=�gT�QZ�z����CQ}@���FA��5��7L
x�M��,Ӌ�}��
��y9�oM�͊[W1�M��Xt J��z�Mb�D�Нb��w�|��+�����[ZM</&��9��K[�ﬕi�k�3�@�<ϟ�������t{�v�� 8ޙ&�&��'.X�E���X�..�,\�������C�RF
���.���JT�����_K��Efa�vn��]�Y&	�<�TP��*��o�2�䚲[ۧ
�4ez2����׎���c��-9ju��.Ksr�n��	��O�X~ֿ�]���5���Q\�_Z<)��C��M�5׎>�������T���\PpMҽ>�, �����n����= �{&�3ms��i���ީ�����P�1>�Y����=�Y3Wa:;7��j�
& � 9��۽��@��0�7e��|�-ߥ4!��z܄�˥G��%&��k]���6Ƈf��9�-ebK㖶D~i�.&��</��.�b�1Eag��^�<����&i=W]���)�z��SC��F*L��9V�CQ��5e��3��^^l�����CB��b2���A��q��Y���hť�3Z3���$Ҋ��EӔm��TKw��G�U[_���h�?< E����OMT�=a�{�ލ4e���Φ�����*��79~'�ɾ�u�uw�"gZ~��g�kVS��y~����J�	�i½�9g�l%�-�]6_��#���24��-&*M�*�~��vrۮ{!�kv�(�V'�t
j�&f	���T�����Jƺ(��20��1_";e#��<��ӶL�̎�$����pՑ�R5���	�˂D���,v�4��Y+eoD�%�?]}�����{�z�<�%n�@��6��_YY��O��6��9�]��He�������f����������~[��_�J�	F�e��ʂ�����u@�{�3�J�T�M<��c����
������.���ELQŎ�W'��F��E�➃���E�ye����ޓ#����ː4k���?��!�>�Cv��.xk�����(k�O�=�7'E��
��8:��mV���0���,��ty.�TX�������ڰ��.Ὧ�z�V3������1�axU%	&�ጴ;:�I��+�q���dv���,���x⃪z��;�xFT���8 JT������ǞQs*�/��q���bh��;��r��k7-hЄ*�}w*
Q�Y�i���\�<�.���{�nk	�G�D�a��y��7��g!Ce��'�׍�2������J`�;,�}�P��.Z�=�����gz�#$P��o�;��^�;z?Ú"�ȉ�����8��j����㘥��,ˋ��{�O��𬋛�n�|����I�w��1K1�����,�{��4�ǧ/)Ws��7��[%����H6��{~�H����6��y�~�$�-%�l+녧�*�j�y�����uܻA6&��<Έn ��Nr~Ì��f��};����-�P��s2�04�0N�V���#e�6��G�ͺ��T�R��@��%5������4� �����$����!ͫ�����	���^7�-֖�������x� Dns�,�Q���[�HF��
_>/X���wR[�,e����t�S�ە)[!���j���<����,v*�8x�?�S^����m��]dRz<�0��-M�xV���}9,7q�~���� �X�!"��y�i��!�[^��'R�KT�N�	��r��%Z��TIyM��7~����e�ۛ���>n��+��5�p������2	a�����-�wN7��x�c��N�J.�|r�>)`M�ů���~i#U�Ej�Xׁ�󹂦�^����<i���E�o8`�2��S��d��O10�r�5��)��2æZo+��DŞ4T�w=��2J��Z��qh"���lJ�6����`�U2��q�Z�nT�ө����-���(O����~�ѧ�u���U�JaM�V�F��]=F��F��8��(7���3��g�K���̴;ߦ�.����L{d�'�R՜k��߹�ۿ���:��ƺ��_/ݤP�~t`�B��ǉ��tغ�9q�[h>yg�����z��L�`�ۿ���xo�~��)��tn�A����~�)a��ӕ��	wC��ߕQ�ǆj3�g��g������rԻ��/�4R���]rG[�{'��`�o�V��w魮��P��}����e���ϳ�*�\�oORW[G/��c?B4_e���]��;����rO+�Y*����DU��O���i���v8��<�\{�w�oFԚ�]����KƪQ(��p�6�@��fi��բ�gR{;�˥ Ih�������wu�������&A�bw[*E?~Ȕ��:�,�����l�ٛ��)7�oc�ﳨ����v*�8a��)�9aI%���?>�(qv?�|[Ԃfάk�aJ�[����~�cN�.�p��j��۫g�N?d.�a��B�*kYL�n6�9�(j5���_(�*MJ�� @w�i����,��Z�C��G��	��H�N�#Dab�g?J�,⯱�������n��ߎ��kԬ�Vq�����y~��U]<�8��qh�m�CQ M�3/(FG/�"�E�����C���޾j��`^���n��.��Eo#�	Zs�����~݁!q%.sG�+�; ��|S��������)��������L/SȒ�zF5{\��{(�i$5sT����ϰ ���F�K�_�t�����y󅦁�b	ϛY�{?��:{Rk�Pl�
x$�P���Pԣ^q۪2($K��d�]���H�"KBrr�Y�(������g�M�h|����&��N?m�����r��Q$���,<t ��dri��j�2H=P�\.���p�F�C��QLa3�*�q�����d��h +�3��^�y�r1l_��V{<�{X�����_�e����b7D�i���J��-�ꎌ_Zyف_�����Ny�"�u�8#J���T�����P���A��m�[��At�i6� 5����hV�>+_��d��TV�ta�3��l�
w�i<;���7В���v�@�lP�ca![������Pԭ�UY���G�9�zF�~�6��w����MCS&�̢ÖC�v��-�
�q��_���a�c���;$u2YP- OA��q^)Y�a���~��/�$F�^*�fNW�Թ��yL��`������gy[�7���b�|DJVwĥ��)����j�Q<MuJ5�l�R#�:%�6���˩ʦy��N��� ���~PL��� ���{qr%V�ty�D��N0י���233�i��7�R4����L���vb�I�Ǌ� �Xی4�=Lq��SZi}$c�'Z�9jc�I%̃g&���΁��tM1�v���RwB~-�xWw���]9��$�l��W���1>|m�r�6$z���c�q��!��m������Lԝ���	�s0�Aj;�
���o7�ĕ ԒGj*8ǵ�Y�xN|ʧ�4�P$ A�?�&Q�S��i�GT�5Zנ���r�h`�3�`�Xڱ�;hm�.��B���������j�U�_���?����SG,��vvz�Y�E7�%~�\�W���*�a��x�%
��=�e�E��˦҇6�Ň�ch����w��+�o�k@d��T�(1�!�F��ơ�����eM�}/�x���)ۧ�}ȣ�4�`�3M�U�Qȷ�̼���/0���e���|��bs�G
�Ozc��cʏ)T$䋕u͜qs�}����8[��nb��ܴ	���⾨���ۻ�l�R�=N���gq�R�o��/���'YrRD&�� �@���>y�4��(u�l�Ѕ�t`%�y��P��@�@
��x5�-\�?�:������>��հ׺G~��z;�_��QM}�]c��C�����������H�tK#%�%�)Jw#� - �HIIw��t	�P�C��9���/��}w��r��gf���~��9��xA��q*~�c�;�nVa#����j�M7^ͺf�3�>�|�)-
��}��#�[���9�)����<c�J����R1Y�rT]fr8ȈI��W��(�=��hHIK[j#��HO̤��������á�����ѹ.��_w�3�ԉ�;E��d�5��qw(�h��4z������_�	;�� 1xG��k=�H��']�G{�ښ_��a�;����֥g@��t!�'�s~Z�&�,/%�;ߘ  �y&�gN����V���3.�
����h�B�V�����{8��a ���&���7��
W��e��k��;}����nJ$����d�x]�z�T���߂�|�����t�Uhc]��#����!BLC���5�b�s��:,n7�b�
8��J��K$��U��G��Y���m��o�ϻ�srp��9��C��=,�1nC��W����aþe߹3g����~�h�������ɛl��O�}�[	x�W%y�4�J�D;hƆ�0�Ϗ ��/�v$����$�����9��贁g�4����v���`�������f1��"��#/�L}�Sax��έ�+KK�m�sk��є�"�N#N��5;�v�
s��szgL�^�(�l�В�}�dlde"P�hl��R����'Y���;m����'{׉S�|��@�3�f�]+V"��l��!�`�ި��-��6��؍�։U;�By�Uc �3Ky���<�w��������W6�M��C+g��w�M��o�����#đ8x�P9"��P�W��L�É��+���Z�����o�#����b$�!S�L�Y㤁:��=�y�dO�N�+�jmqmw�r�� ���r���V=3`)�ؤ�3S�e\�X���,k<=�+��
\HMD���^nx��ާ����gO�p��D��h,�?x	�-�O�(ӭ��Fl�<�Ck�e>�Eg_	��e�S,�E>g��D�
*��[����pEy%�JG~�
*�2L%��;ڟ� V�CgFd���l�Z�>�c�&��-�T����8�T�$;�(иs��Q���7KK�[��h�M�{�
�hl��!z/��.���2��Vtfn��IC( 3�,͛������O^��n$�c6�� *6���������U��k��r�#rک>J�]�>�����b%�yK++0O�x�C�;��S;�6 v��|�J�?H̿o�x>���mi��q<{�;1+<K�"Z������^:-�q;|1+���j�����+����\C�dGQ��Uζ��ӵ�<�ZN>�$��og��"�~ڋ&��Jc�y�g�g���
�L����ʰc�{�7'��-Խ:S�:F�C�%���V�o8.n�5$v7�uZL�3������k�����8�|��733������tW���P�%)(��o���Zʒ�λ��ٌt[m���n�=�ZW��10�&R�Y}�a�jA��Ӹ�0�1y~�N�
�۰o~ ֧1��=����@�!"c���mc����G�.����Kg)���鬮���&A�Xs�R��f�O�s@[�4����wh�_�ȴ�uձf
P�H��(J���z�f�k$(����<8<��Y98� �6�\����c���	C��C���!���i��_�"~�%py��s@�[��G��
�}����8����'�u�O�(
]&��`��h[��+�;��uO ��DD���H.��w�"5=�
P���؜���e:��K�\U0C�.'�F21&ڠ�Jw3lf�ݦ��:e�N�������D8S��;���D�(m��@����xؚ(��\���#s@�͍�DK7���N#^�B���H XA*�ٗ0����%�������� '3�	4������� DX���#��7�W� Z��Y[N�I}/��u<�E	3�Wk���|�Qic�Lx�B,Kt�2N�]����`K�쿹)80D6 Wz��Z����;�����h�Fɴ�Ƿꞔ��LU�E���Ȕ1`���2@�[�����s����vfV�����u�`b>deQx/1�0��P�Qh'�-��,\6��/�텓�LC�j��Y� ��	�yW=�hϗE+��1RRR����s��e�z����%RG m���Y�6"�h��%�w����jq`` ��=����.�]�����1dLҸPaξi�d�<R|#?��C� J}�'%��[S�̺5z����yMؓQ��2��kdf*����M,�[n�w��!h5Ba��,Y�n~���EӬϹ�Ҿ;]g�9g�>`D&d�|l�B����Gd�W"�;V���OSӸޥ[Ih"9�]c���@QFk����W���t����9{N"�=i�q~���/-a���t)���[��� ������V���w�������I䂹��*��'!*������;(��U�Yz[8�'�#j5�K���Oc�ܹs���-C�[������f�}%�a���D{�=qő��L����A��L6�Q�Qb:rcI�#;��Ye�sq�==��7;��ҷc����_�d�:�id�,�1z9�e�9���!������r�K��N�ʐֆ}Q���s��m�OG���!��;l/oo�������� b�rP��=ز��U:5�P_V���� ���Z��$�y��"@*��P�͝�ƀ�f#�v�׀��������˧��GT�+�r��zL׮9W��Jf�ѭ�[��y�	=9�z�EJ�J�g���jz}�E˘؋���O
D��<�*�o*����-����Kl1�w��nNHA^�i����獭#���{�d3�tI�om�
�nYmMU?h ����W찈�:�%H�E��7CԐ�]�@�X���@GC[�Q��Қ���������R����p�>���֑��h�e-��,^t:R���
�%~H�����I1O������zQ������_��{��ť��פ��[�bF�K��:k�|!{0N�yW�� ��_3Ύj��2�U�W�ˍ�ww2P=ަ ƒՍ��Yk����H�هd�k��}]p�QeIDu�R���������$!!IIJ��������ZH��>o$�n�4�ΨaMFH8��$��!��k�㓮�ׁ��9[7���Ҋ"@`��&Pz�r"�=ߨͥGRן4�����M�V_
kk5��X��<}-B�\����K0�`��tO��c��T��a^x�W���]�r0eUF��O6fye���� L:!���Jˇ
0�yW��7�C��UKݗ]�\#����z�6�]aR9��f��C-��q=��2g�Z^vEƗ��<�����~6744��n8ZT��0w�䞞��1;���v�P��ǳx����Aن��������ihm�[��C4�!pf���r��Ƹ���;%����@;[?)�������l�D�gz��e�Z$�� ����d�Jr^!@L��ƛk��˔<�,�5�	���+岦�a^�kѣ� [�1��P�Js��1��"2 �WqR��`��̟�e`��ow$�΂c i22nf�I�~=P���4�2�z�~*(wdo�������&��J��D(�\?|��A��S��jA���{

����A��.�ߓ3��lc��8��������=$TB<6�!����A먶����x���4DGGǘ�NQ="�G5�#�9ZL���@���°�#TTTB��^o\�u���R ��Ϝ5/0Ho��lN�}���v
�4�1춎>��@l�%�7���/��R4/%�ۥFVx-��qN����ùh`_@AA �cI�B�	DP5��U��+C�xg�R�$ײS�¯l
h%�*� �ڐ4�� ��6&���ނK��Gn�����<o	f����qU���=pam\/��e\�/[x-�VĜ_/���� �MO��<�].�q�p6
�Ӈ��9p>vZ��N0" 20�G� ��~�Qw��p;WL�b>H>���_�6=ƪ]�$Ϟ�#��Vh�Aܪ#�%�8<~Kt�,�t7���夤��&0��Jp��}&�x
��P�ܥ�v��f���*��0�F����yˬ׾���ӷ��j A�ٳG��=�!�\ 	�r�:�icIc+��9�~q�t�kp!�3!H O�O��7�}%���?�����6{\�ϕ�mbd�x����2�N��4�`���^�ƣ�y��<�A��A�G���2]ƙq�q*��OX�i`���Q���/e57$����
�7��GGG�j�'���MsU齏��6�ZK1}O:tZ}�?d�
l�D
��r�|��G2$/4O�
��O��#/�2���MMiT2�������0�@42�b�8���r���֮�0���|lb�Qo��ف���nG�V��5��H__;�x��Ӗ��D��O3ė����>�&��T�\�|����t�taB��7N�ԓ���nٱ26�XXX��}<<<�[�v��^�Fؚ����7�m��~9l(����"5�)hg��.�G�Z[�0ܾq���c�p��ȍ�;o�i
�yy�\j��"�~���ҽ���f5����Lz�e��Wz�O[�vD���d�8��~�ꒃ��q

꯱A�d��8��3` #��TٓGݏ���*�B?�d���2w�ϥ��nb����bn���[Pyp����~`��@�ǟ�Q�8�яQd���n''���������<��;����#�BDܲ���uZ?�88rV2|�#�����yy�� bC6��Ah�Q7˄�bE�����9�Lש����|�n���M5U�C�+zxx(�󰡱��r��(��[E����S�?�p��fJ���Gvw?�9�JK��:�z@��I�����;^��٫!���Jd�&-Lman�T\\jn�����êh�)y^s� ��^[���YÅX����zY[���+�yGtӫWZ��œ�R�	\������8~x�
���e�Օ��������/�+Q�Z۱tAO��F6�56�t��I^%�\�Iڃ%y���D��h*i���}�.�e����PSC���:���=dz Q6����*� tK���s>���HR���@M��N;��c`%j:�c���Xnƈ�>����#��z--�I��� �;��*b��2�'�#�R$��-����������x�]�
�1��+��>[��m>�-�߮�9p����h�-�ڭ��,�FW���d྄�&���i�P�b���(�����̻P��7$)6��>c�� ��@=�e��U���� v���,|��ݴ��5��x�šP��[���aK���
��!��^���c�>Jb��CK�
шߔ���H��î7��bM��� ]���ͤR���w��V��s�����:�������+�_/����-���� ����"��=�-d�A���P1��~���Gl�7���6�xg����/�`A���H����ɱ��ފE�H� A�=m�ݰ��Rp�&�UcS_�8���nЖ�n9��au�m�!�k .^�����_J���QVUN�1
.<vh7�o���Es�WYѥ��@y,� �a�E�'9`$)�O[ʀ��ή�[�@O��=�U����^`Ą�8T�uЕ��|uO��ؚk5�k9���V^^TL*'e#��a�5���Apǿ	�Oa��������5!^ޤ��">���t�t�pxo�A��3nV@ՠw�FF�x�%��;�u����Of���11����������2�7�GQ�d�G�C��U������+T��|�+/^����XZX@G/�N�6���	�.�z,'���:��EJ�7����$�z,��BC�A8<?���K3pH�9O�Ș��#	 �T�����Pۼ�VU`֘n��SeR<��ص좏zL�����������2���daz:�21@2Y��a�. pF���ƝsG��&�z߄��<NKC-����?k�^^M���M`J8�<��C_�M}?Z���+D:7�!�<����)ͱ�|C)�G\� Q�ߨa5^m���=M6� 2�c���rr��K	�_�{���;Y[�)ݶt�fYZ����gC	@'[9;4�4�� C�xyy�d�ͅ�Y������j��&B�r�:�%}�A�)��bG���R��/]RR����cL�jgg7�e~cֹ�J"v��J�Jچ�߼��V'H	�Ywi &G
�����'���e���y-���0(��wa�4�%���q��/4�8x��(HlO��7��#P�����s܋H��y��&���b�k�T�{%e�ӵ��M�sw�&��,��Ӕr��ąn]$ ,��ĵ}������R�ٳg�L+��п=F��-����n(@u�������d���]�ѸE�⩇��=�>���2@�Th�x�� ��:I��RF��,�X;���2�n;Pr%���.��wQ�.ll���J#j��)����y
,T��R:�?^��/�4 q s=@����%(Xbs��E"?���V��9Z�Fu�����Y�3��9�ctK/G!(���3��he�𒖖���#��׻tt^��ns���]Vb��T����KD,���ܪnn��C%��J7,��~��I�������2��ƿFio�X�V��oK�L�l&y�����C���g&��xy݇vD������i�l�A�&Z�2~,���� ����P����񳖺�^bku+���_9�VP�|$�-m����>��M�ޯ5㸍�f	��䏛�nF�}�)/@ό�E���$$$�VV�6�4��ٵuff����m��P��m=;;�r��1��,���ЧC)������Ȥ�� C�]�������Jo������&{2��Vxxx�)=,/��8%�IO����k�ptMeL}��f�gK�?Sq#���4�������§y%�hN66����ԣ�>O�꠴��ܳ�ć��s���g�`�lo�܌�pu�����s�<Z�-�V̇P��`��|����weeZ�i��q��g�^���B-S�,L��3i�_����#N\Pb�˖����	(��8��_~����*�,c�6)J���p��� �1�y�gg��3�ffߝ~��������؜:�������22XI�?y��j���ۍ���ө wX=�3�'`�GS�*��!	`���#��&�B��c���)�Ig�N�?(|��|�U&��,�} ��)���w�@߁b��@�X_[JᲒ�����?�*��h���9:��{�uq+�{r���>Q����BzE��������^���\U��@_�����n������{�M���y5j��8�+P�Q������@� �<��g�d1x$P�$���=xP0(��)�B_����VQ*���&
��榚��{]ݱ��Қ��ax��w�;G��"��^hm�ƫ��4u���y8=.�,m,�2_�������*���[Q��w�\��P�����VNBD���� �2Kn��]��_��U��>�F����6�E��p��i�e�EJX���|aikz����Ďì�{2ǃ��W��O�kk�����^�)(( ^Vur�|Q�P����� r��4��7cv��]�4E�?��&h�aL쥏�^3ζ�!�ݛ�m=\���Pu�qY����xJ �*�<V�N��E����HEق��f��$�{��\q+!_����*�*�����(�Rr��g�zJ�#��#�$$͋�:	��K�T�O-hN�9�nn�&^SEw#�ofdy	���
��ڝz�t��nL>X�O�E�i���6S�~���1�i��Nrڨ˹E&Ũ�_� ߀K�j�����a�<��_�6y�[bE-�!��K���*-9򂂗�B�{�τ@�����uK����\27�߷���:�2��PHH�6���S��־����G�������P�=K8���7)�����O�^Q[�ݟpI���k$HЬ�ڲ4��F�8Y>M�A���Q3��K�à���6����K���� ���%�� ����g-{����'��)��-X��3��)�W��߽>9��^�Oo����މM���z��q+<K0�9��7����3�^ٍp�0w�*���{F.��ι������ﾃ��� �/�d�c
h'ܐ̵�����s�S`��5��twx~����0M��c����!he^Fu��P.��G�ed�.� �o��r��Pu(eV$��g���4˵�ʵ�">W0A�cxxg��Qu�_��0sr���;��L�E&�b�?5IFD�-��]x��"rI�e�L�����겇���!�\�T7���HNo��o'�b>�APD��x�'������C
��w����O2M0���O�����b�2��Xߵ� ��F ��� ˈ^�퇍���LR&�[)h"c�p�l�:��5����K��ؗ$^���R�׬4`vh�� �z)"cpZ�{�T�\˺3l���
�(��X,B��o7p���7E,ۀd�e�Gl�X�M�Đ�A\nB��a�d���4����I{S�`C��]���(&kJ�y��-��Jk�����,DQ���Z�--��w���h��H���,Ӄ Rl�ЂG��6�³ #����Ng��axI��Z���N3�n����#	��F�8b����\�p���E:(o.*V��L��t��G�
}��zG���i )�A�W7=�r�0h�H�k`�x�噥"YO_�[ )d�۔n�(��S9"�ɁLhY�fYM���9��<jʔ�>g��/��˦>��'�U�K�d�S�\�8�ʰ~.-%�D���!���\=���[ )���
�����^��>�����v�?�tz��8j�Yv�id4��*oʃ���?����s�[���2xJ�/�P*�����θy�͌�]X���������;ؒ��6%jŘ�p׵Z��|�:�9���=h��'o���������κE�l������TU6.f����^щr=�ˋx�&I	�y	x�fR8/J��{�k�5��Jì�C�#��IVƔ���w��%�bc��
y�K�fӂ��I�[��ٓ�+ʌ�dnQ0��T���� ~n]��y͸f�]b�F��nuuI�e�8K͸>6#��]~jc*���c��92l����﹎w���I��&�ȯ�����n��,�E1��k{F�))� A���K?��,�PJ>��.��Q�����&@U;9��y`������1�gx.�[���ǺR���-]qz���ԁ��ԙ�欪�P��C�N�L�]���]
B޴qAte�T�XҺ��c�CN�t�&����Ƶ0����:������g���ɂ���8�E����T�j�*=�u;�R+9$$HΕ@0��+�HH�IB���Թ֚����@�c�/2�_}O�^�s:${���h(^Bۇ����||N���� �Y�ԯ��Ȝ�I�;��_�%w7잒�}�z8�?�'DE�+_,+j��2%��Q�s���Z�j��-�C�:&��ȱ��.��5J-�in��ʢ�)�'�w����P�X��R�	�}zd�Uզ�5>���+�Vѻ�c�x��;e�˼Lr�G%�,�Aᳬ�ni-���������j珘n����=1>D�{R%�4f�1�5��K�ϳj�v��|RE��Û�lB�tsS�y����j�����W.���/6��cN���Y�GK�E�;f�i�/#B6]����n������v��Q	�ѿ}�"��l}��6��A�P��H��ZJs��H�V_���l$^-��?��X��W��t�|w@�75�nFV��ωԛg|�j�`@Q$��%,&=$l$t�����S�(��u�`4]d�&�'d�G�o����q�?>�
��_TSx��g��:��=�mRp1����^D�U*����_�ñ�oM}����ΆQ6��2�����}� C0�+o�r�}NG��4m=}ve�^R����w�w�v��o}�����i����Y�X�MJ�Y;1P8��EJ���c�jsN�5���eNB�ߌm0|+�ۻ$������8�͓�?�N׻��\� �L�;��0�c���,��(�S��p|�ʜ���5`{DR��2��kԜsвZ�!~p͙t���N����'M���-'?��jrz\���D��6�����Q�����%>�]~nl$ZMM���ڹ�Th��1���p%	"�V=V���=
�,��e��0?����_~ԗ+lp�ʴ�O�O:%���Йoz�C������g��HG��)f?OuĦ4-�X63"�$� h�?!]���^�HM�FQ�m��׈e����/,`��D���KHJR��J�`�	@�]ZR��o����xz����������IvV�i��D�[����s��m�{ٴh��\!ݺ袹s�Cn��Um�sL�����+ � .//_!e�!@��&8�Ü3]w�C�ϣ43��H ����N�KHD���^ZZ�r�e���|��Q�oT���(ŅWI��kX,a&T,���&�W>�9�~�V�|�-�=44.nm�4??���rWBJ�9���5?h˴���֖���(�k��DDD��u�&�𖉡��T���*Nܟ���N�\1�<I����"����q-�r�N��p��5�;�ql2J�[O���UU�����~� 9P�%Y)g�\H�too���D��o����Nd\\\�<��B��;R�t͡�u����}�~I���z�KP|씠d(�aƚ���#$*̒�v��C^%�޴�V�q�]���9CwaI<���Q�W�X��eV77%@l����w����t�����#��8ݟ���L� �o�K^��|I	��m���6"s�>��.!�M����fRhh��R��(���x�Q��;�?n{�����p �Zfyl|<;/�N||��u����j��"�/z�*��}�)��ەr�Ya;�!JF����Y�1�Z�]��iM|�p[T�ٙ3&&�]zz$*>9;�#n�G�A��������������Ȋ
���Ĝ�\��].�^�웟.���Tb5^�a�B˥��F����{��|�Pי��ꇉ�
ntj��P�G�TT�`� KX�ß{xxd�Y"�>I��,��M}ਯ�oEHGG�+��72P�F��(F�.�/3���QZ�aqͲ������J�wd��ۜ�R|�V>���wycccr

�����%��)s�+M��ss�@��>�W~�Q;�E��H�.�e3������r�:�q��ylE�ō#ﰣ3>�A��D��*N�4���{ڄ:�ث�U�RR�===`>��r`ή���{<Zi̙���ܛ��EFb�
�����&=س>�����Tޟ�a��U�`&h�Xr6LI"*�y����Z�s�]���F���Opg�UL��C+�?�N��:��+|�q��$�"alL�<�u�"s?��{Cè��;���hWa��C�����>6���ڊ]��(w}�8��du�7�fV�O|Jg!g���qtt|����iF��Q�:,4TT^�t �I����^���M1] tyyY����Vl�S){���QRl�h��b|iz��Y�t��d�C|���1u�.=9[�Q��{���8,|���}�\4F�")!�|g�9I���)r\w����1����z
ۇr�V)�451-(N�Ho��e�kb%��K���DO�-Ĝ�xLz��׈���SE�����&����5F��j�u=������`"	&���9�f���rr����3��M��M�<��e��o~��>�� ���~�E�w�	s������+vVY��KN~��_���wqᵸ���:��;���q񮬬,��0R���C�|� >�y��r9; |7�Vo��$S$I�LPK�T�5�k-�� v��!���9@/��1�x.HsKK�g��M��jk����,,�2����3̼x�)����ɘ��d��N���m/�,����@�a���rww��Z��R���ۏ���g|�~�6���H�b����� �����[���8|�χq�J�|���S�s	<=����T�Y�dR�((���[ɥ�n��fgf�F򕤍�?<xv'1)��ɰ��7�����
6
*����C�J|���ũ`�k��W1-G�Qz!Yśaˡ�����Ŋ���K�̽���U�g>�������S��Z��_2���m�@�k���	cv��
��Ǡn+�����,.��?����>�mT9����2<İ=��;ra�jkr�wH�DK���ˀ�(���or<6�'^\\ɺ{U��4�Mz:)(ٞK'|i��
�?�����?;XM�id<�3����~����~k;�s�Se��λ���`t44H��$��$;;�)��H!&�\�DI++F(<ZZ!�|���&��{���M���{�bI���~�f�vv�j;�T��G���5�_�C�n]��to���$�l���_⣐��V��1�Z�Wg�����G��ض��U*o���
�����oj�Ѕ.�m�k1g�M�ؖ\hT"w�<ƪ�xr�!"J'B�,{y�8�q>\t�l�Kh������1����Hb��j�s�±u�9�bFe=��55���T�$�W&��e3S�{r�5��a+�����N	>@T�t�Stl�B�s3�h�z��X�﫩��Q�42��t�l=��t�^t��k��I��p�,����}�G_)��(b(�Ia�����+�+�iʞf5�&�� ���+ʅ�?Q�v��سS>>&k��|�~�M�Bmmm�P<�Vv���H�we��L'��~���s�W܊B�?�S�"
|�l�İ4���Ո(x�$���e�aw;m훰��������h̚��'���EH�����>ɗ/�"Ʉ#����\v
��KW��:BR�g�CC����F//��/P�1KOcb��z_�k��)�q���R03�k�9 m����ݲ�˯W.*���3� ��B�+�z4/`C^����}� Gh��Ej����ݓ�i�?,x�����)���D"���£�?B�Ȉ�H)����e)P��|�w�d���J��i�GB�����D���4:&&�Ouk�#saA�d��y]ؼ���(�5A��-W�����宮���p֯��Nb-��zz�� _�]]T@Q:��w��>r�8q�a]�r<�&�������P����`��+)���p��� �4'
o�������r�SG���
ç�|$	,�a4r	�uu�n�_@��8޷�iL3�=%�:j
{S='��N��PHQA�@���6���?i��������'�~��D����~K�fR�ؓ�%&C� K��\�h`���P�l�ԛ����b���P�or�G���	�̬�y�H��U���s�+!�gӾS7�9�J~n����%:::?�0�����܁h��t����G(O�}���hr4���N�q�N+����u9
r�N3���kp^l��^o`?���.K�Uc`s��+֩FED���k�ۀ-�=B{��|l���O�6p�PB+�	���I���=�GEy��<b��x��T��$��^� �!v�Y��iA�ѫCQN�]�n�	?�����6S��I��Y�-�������;ý}�E��Ǳ*��c5Q�Y�߸ێL�V'� =����5�"���`>���Ob�9]��\>�,*Z�ɗO��cm�]�:�kSQW�S^:��Sc�~�>`*�Çے�����G�	��9{�z��Y�BM�Dw��9t=��s�_�!"C��a?�i��D���ZB�k�i���R�}�m�����J�Ԅ��5��[���$0����~G\�e8���0�(1��R�0��쑉K��> n(f��}�=g����CC������-�r��������;,̍Đ"1���?�r�)_�r젓�����~m�׋�Ť�e�	�1H����~�òCRS��S8�uE�u� �{7�m��oT�\I�;!F�Y>�aV��ĝ��`���问�Ej���5{h�b��5��%%�0��@G��(���{}���S:��'~�͎b-,��UL��}�Y��_���n�����?̼��J�!~�!
��DV(�л��\�;|���"��(�����nZZ��i���H�YzYʐ�z�*��'NBt �?�Q���n:�}c�_��~��ƌ9��޾�Ty����Q�y��=��<�o�]�
xhP�O�oC=tϗ�~N����/.�CBC�T>����~߷�X�L$��"zNNN�Q�,N8:B���|o�X_��ج:Ռ�U�^�tP��Jďϱ݊�t��K�R�
������	�ne���x	��R�үY����2Z�lht����� �ɽ�
AHC���*�(0Y+Jo�!u2�0>�_J�a<(�͛5,�	%���.���;ctg>$A�'��UnZ^齆1iOt���Asp��K��q,�`�����T�m�{}j�)̜`L�f���-�=n��n7�.���j�֏��*�����9��
�YrA� ��֣�}��}�����]�8?����c�/��%O��#;�1��k�gt?!�`�EP�k�g$��f$9���h����'S-A�N˷�ẑ����Q���r��3K&''O.�T���ܳ�r�W�V���w?��&��k;H��67������M�Л�o�wo�t�p�NV����i�{NL�`�S�D�fa�s���k���^�,'��v���M��uT��HJ��L��ۙv	�P��𯫜����n!��Bmj$pB�O��鲛�����^��� �UwyWQU���sqq!]�o�;���A���ХCR��%0�Eu�>�^�;�6��HS�H�7���S�e|r�����s� �
JK�n�4���5��������z�����=�o;�,�*C���+��'���>�@�y�E6ѳ�b������^�o�i�{���-YW�˼9{6,��բ���4n�<�	����a�w�P^ٜH���v���w	-spq���g��Rt����x.
����bï�������H�Z��S�f��gcHoƘ�?GNM���r�>!Y�R���]{�.�������d�Q��ɀ����U+��u���oAÔ����1s[�ga�p��;��?)3���(X#�E�Xb�52��r��'T���T*6����v�#ԼΣw+^T�ߑ�o��N)��Y:��r|D�����*䴟�(}4l@����p�$����Y�Le:�$�ņ��_�<�E�$4�t�(���0���X����*ue��K����R���#���W$�V��<����tku������x�-�^H����Cl�\+W�h�ɝ@�G�uk*h���;x��=U��z��+,���-#g���\�J��{{zځ����Y�1^�u�n�+Q��/���߽斖�y�l�6VKOn-�6�}�s�J�	�7�M�����k�wK����Iv+"�������=t���-7at���d�%W�]TԎ����c�_���m̵��ב�o���օy>۽-�[z���֩i�z}\IH�`
���n����#�α5Q��`=�n;X�8�Ǳ���|/,����s���A�r�	ޠ|Z�W�j�1~�!��f�M�vC��5к@��[�1�d���O�WZX�|�����;52�_wH���CS�o�S�5 ����|a!��Hr�w�>�
���u䷕4-�v0l�\���~sNª��O\򧧧I��<����:��8knw��H-o��S��G��wO,i�m"<�>�s�/#+�y��}tz�v�s�/K��{�񲸸���� a�f��lc��ϵ�|���cy��q�F@L�J+��!�(��>����B��P�S���`�̬����%�C9����Ƴg�pϞ
S�d?��u쎇�5�6R�����*������� /qpۍ�- �Xئc�Y��A��e�JјV�+6v��\P��1j����`bv)pϼy�a�s)��Hk�Y{J��R.�k	3�n�`������f�zL�x|\'���&�\� �f�ߠ��-�)�N��A�~�kVC����'I�o.���Ѝ���79E���Lq�ǁ 7�ֱ����_86bGQ�����|o��
��u�w��B����9��JF�����8	\�oD����
Z�F�f｟Y�!���a�L{���e�7�,?HX|����}�B"o��*뢐�Hhϡ���˗`ʃ��Shc�uvvv����e&ddD�}�&p}�O�̼��"g-�h};"߯I��>����!238}B8w���$O�c[��q=�=�Q�2�tJ(��Mȁ�H���V�Һ��1�XDh	@�ORv�?�`"	*�e���+���-�G����#��
�E7X�Ơ���-}x�I:��&�����	^� �ң���]Lȭ48s�L�ߊ@H��p��= �\1��sQ�	��V)�/Q�U�i����BDW���.T�]6�EW��"��~#��4/����k�wy��wZL@�hs<''�u��n-C�20 /����}X�q��)��bf���>*`�r��9s-��_8K�]x��Y}�Y<((�d^X�ؑv���6`��]���4�sK�uZ�L���9��u0�@�EAJ`��w�_�?.�1�����*��[:�s-$R9C��)<{?��5Iw�H~9�Ld�t���u9���܎n����VR�R>Pz�һEo���s_��^wSt�|��pͤU�y����.$2.rrWy4Z��� ������ZQ?��������d��[�v�U��w~Y��ꞷ�ͽo,�f�?ź��'x�����?j���(Qq��bO�G�$��j���3M��yw�~���i-������)�(��,h9�E|�L?���P��zd O�*~��齅�K�.�F8��8t��e�PX'����d�T�)�����gi>�v�/��C��jU[���Π�)�8(�g'����))J��%L��K�
ls>�e�{��4Ү���r��;_:;Oy��W=6�slba=Ɵ��N�W<��@A D3t0T���|�/�%*��9n��C+��}<���uΣm_TX���Ə"��E/��l������C���g��B{l�WύZ�ba����� T]��C����48��Α�eϲ�"wsG1c2�t�?���J�K���Ç�3.��B+�FFFEE�no�e�o
�k�ó�邳KhK��4�'�<*G'&���HV�:,~�M	�7Q�H���	z��}}�ax��j���,���
�-��؇e6;V<�ݖu%$�]�*_�Љ�/'�ϫ8�����g=�W�g�B��X%�fd�Q� 
��������V��k�s�@�k5{p�ZVc�"a䪆��<�z�����HX���д<p|��D��U���_�[�q���=?�
�6JĲv�~�����1�m�� ��\-`�^n]{����z먪��_���8t�N��D���;�	E��� ���%�������{���d8{�91�\k�H��d�6SR�;'ȅ��P�5?���/"�t�+��eRg��]o�g:��Qi���;d((��R}�c՞gf�s��/��F��ӷvv6W�c������ζ�nj��	�]�i��h(�xS�'�	�����z<���"f���rbb�q��㢌���t�A�M)}}��"cc�S����6-��#"m*[�)��/oz,�e Qc"~�O����h�^���Dn"��+ �O<T���100|3X�������
�^���x����EYpa����Rr�l�\A��<���l��j���a,�(�"�t��ܟn�$4,��Ċ**G�0�腋�dߊ�����at�ׯ_�r�᎑{(����a��i+e���ݍwFB�V����]�w��8� ��EԋU^���n�� ���a�O^�qb8u]�����\���'�N�+v�H��mfL|�����n�;s0aO���Z�D;c�k�����d���'��q�j������r�8w�%/���r����P�J1����g߿��O��z�Ժ��'vc�w�@7�qǭu��ohh�a����	����������PI��t��%�������]ZIC?�MQ�9Q�|�}#<����>j������q���� �_n_O�iVW��:�?ߗ%���$\r���|���$%�)��/r��)�`�w��#4�ū,�~��@�)k# �����wm<�hN��y۩���so���䎌�J|h��z_�xq�|�O����H,
x�W�J�����סEC�_���jk\mr���ui�����W�}�.�Հ,dL7@����-z�@hA=������_��_^�,ں��o~0nxF����;���+Qh))�Z'i,^W\ ��R.Z��ԕ%�|"a�KD�� ����I�r��/0Ub�p`&�s�/үa�����U�ݨ�`�h�~��=$id��K��X 8c)�FW5���;�:��T+lll���ݎh��oF�p&#J�)�unl�y;����!.N�����2�q��=WQ �Y9�1��P$O��U���
�������zw���;�ߜ���<�X���� /l��#'ߥF'�j3d��+r����@�J;;;�c.D�+}��Z�Ϝ� ��'��<��,�[J�K4����S����6$څB���r�����y�9��Cw��y��*wQ���4.phZ�}��4��|�j�o�,|�9_h�0Z��fМ0Z5��-��9O�.��M��}P�*��RS��ø�5;����X�>���$�nc��+�~w�4LF��o�B�=�4˦a���!�%�٢�iNwB2�1���(�H�-Y�'�\���r���`��/19����Du�K����.r�?8�Cb(�<ɶ +	 ���p��u��X�W��ͧhK����������|���-)>~PE��i'j��ye��������u��m��|1u��;������i)�׈/�}�x��6���6��Y덏���������*�P��QI{;�L&=��0�ri3��T~42Z��^KIn��.M��/e��9=j�*�C4���ɝ�X���ӵ��f��8��}=�7���2D\��lm/-Q��F� ����߾�HH!��5'e�R���Ӻ�^ڢ��y�kg���rsss]{9� vi�|����-HJx��#t�R��(ȱR���+��KGo����~�ohV�d}�9ө����IJP��llN�[�aS������jj��;�a��:C���عM.l%.R3?���>�u�Y�h .=l���8O��e�Y(&��5�g�~��	%�U����,�o���IͶ�kE�Ԓ�� o�^��"��`0�X'!��[�П,x�*�id����2���܅p��G���ߨJ��!�p�[�hO��}.jv��Ƈ,n;��#<+��f2;1_2�����	�N�pb��(L������}Y�m�f? 1��V��1�n),�w�WH&�98�1��L
�A55�c:/������^��;> �����<v��@�ߗ5{��1�؁�|Ř$jQ�ޠ�D�G��!����3)��
��lQq*Q���G��h�;{��d:�̈�3���3��s5V��z�(��*�TTS�;jX�/�������L�Y�[px6Ľ>��Ո_�A��d�JBW'�@�_�������D����]vE�ϾO�A`�P���������	���a��d��MŴ��*P�yQ��|��)���Eڧs�P�m�K��}�M���n�B��(LL�
����~G(A�3u�F��NN��?=u<��A�!�|s"	1qx�IE��HOOo���]0������>7�ٲ���Ѯuu���*/j���k�Ȯm5Cd}�׹<٪v��tLL��ғ�gֱ�)����T���TWPZZ:�ĺ(�\�:$W�����)#����A�{���:�_�(��)[�#Z����Omzz{�s�*0��9~�� $HW(:AbN���9�3�Ъ/��ぱ�����0�x����\�H��.��b֑[�%�h��*��/��W
aHt�p����5�> �L̛�����Gǹ.QuW��<Q���պ�O$V����q��n��]�JG���ŗ���"��T��A���BF�7����ҡ�"�HOn�\�j	D)�i~�0ڰ��r���9��w��[��t��/V�fN's���Z�zO#?�U���g%���N���� ��
Q��KCӯ��Zw��������S���K�^yo��J�Ԕ��7��"#מ�t&[��!�+�����_[��Tr�r0����0�Z�Q��g����S��0h��0{R��`�����۷�r$R�E4o2��`�F--����-�(q��'K`�2��a���v�n�җ�P%wO������EO�� �zG�lv�;��d��/�x.V���-��Z���RY�p�ka�BT:���KZ��� F�<�%Rs��U�Ȼ���F["Bm�����|���Pv�;� fL�`�NBd^B���Ng�h��ѥ���	qT�¿�
�����p%d*~��W�e�X����ETT���z#�2��y�¶D=Ry:M�i������ܗj�Ҥ�/i��bTf-NO#�� [,�\?��������\�B�4G-���ѐ� ��O#�K�����̃����ZWY�9`� ����e#���A싧
��=�w�ݪ�7�;8��6�a;t�$K�%u)���lؖ�Y4����ǿ)�s�̓�E��[�sttt�qL�x� B��+'���.��S����'f��#s���g�YL�
'q{{ۯ���a(�5��H�Vm犺�q��n�|��^�����rH�b�z��l�u ����,��$e͵��~�]��m}���|���ɇ��x�	䰄ҳ��3t�nn�pm:�6v(P�
�І3�[7���Y�o|�e�����P�+N�� g��A��*�Vu(�b�A��hBZq(����}EH"o�G:tG>m���j��6�� ����I�����w�I %niJ���=f�t4��
d���$$!���d5�GA�n��"�Һ��M/FG��/�V�D7���:�4Ti�VP��^GwW6����F��"��+�c<lU@^�2���%��\�?�gY�4t�qeєg���=���c#@;��沐Ϗu�B�N��Pq�ũ��]�0�3���AߵX�ߗ��[GGU_�<e�������0��`���ޫ.ّ&����ַ)CP|�罴��XF�1�2d�Ǐ���T���,�L��jg<2��)�I%|Æ"�����!$����H��F�H�[��mXf+�h�b�s:�%����x��1@�N���(<8�۾�������U��0@��A�Z�:���
�q�I=�繁�����'��U;��u�)��������<~s�000�ؼ���;�u�����Z����w�ҺX&�YwVu!P}�2kl^��ɕ��6p
�yV��e{��8R��0�v3�
���d�͏��F�ER�Py�R�to6q�8��{��L��;��Yב��ʊ�����*<��~6���5���+�Z��Ax� @��Fv���\\�
	�G.=�!jx5{�h��jLC��S����$[]�����Z~���8����;���ިYe�)���e2�fA@}�Y���3,�_�ˁ �G�V�O:��r�o�v���ػc�fP��X��D�h�6���E�ѯ�tL�E�4S���7�8�E�F*��K��q/�����3J�T��8��H0�Fbe���FvbL���o�����߾�J�����Ǆ�_x�O�t�|(?\0����\N��l�+�tc|;��Zf�,~�΅���zn�cs����8$����/��v�h�X����H��"���9��f| ��8K��.�u�*�K�g�PV������Fb`�}!�a�fKvtry��F	���l���144��di{$�TK}�2�'��=����B��0���6,p�g>��KGk�f`�R'u�X-��x�>}�*H)��~��!�w7i�����O?����=k*�0�� ��d87���h<�܆F@�6+�up�R�v��0�‎:�	�m��o'��f8�qF	��l_y4>�꽂�t���o�F�Uqa�U6#3<����UGͅ�ƿ��������p�)����Փezz��o�c��~����N�OI^�!8��8ݜ������F47c'MrQ��W�{�_�`,9qg���g���V��Q:w1N������W#0�FFF��m����3��F#�G9��*
 ъհ�uXay�L�Y��s���$S����n�dz��O�aSl��	�}�m7f/���' �,�����w�TY����Ĵ�p��k���	�i��LR��n:}i��s�o�D�d�*�{R�c��O֖蚶��M��Q�͎��D���� $�g)G�~�������{�B��o�~��W��Zl3#q$�Ja24�0�Aa�!R�c�<"���S �*�P-��C��Y��b�V�J%����%�Gb�I���S���/�){#jI����}(3l�+���bR301�����;WOV�NJMOg``�^���r����p����C�я�j᜖�y	���UBi����L�W���qs����3)��M�A�s�v��J��� �-��EN}�*��`e�g~�ޣ�Tz^�i&߃k
�;N��޸���O�<cbwOz��i=��$��|�VU�O �*~�=��wǿS,s���{{��/��32HA��$$P2>�g4�� ^ۏ�e�p&?���O����}�nD�2��3B_e��o5�|��X����O=����jg��T'8�t��Kdx���HM���7`�0a��v��7QE;,!�q�هD��dD>T$P�ľD��L�y����m[-��T=6�됿ӛ��_ZQ$9��F�^���NF{a,J��Ą��I.�E5.~�	��&r_��s&{-�4���2|2t=ɖ8��3�Aڌ�9�����@2�5���8��;��_��<�+q?��!)�E�b����藄��=�Y�|���fJؒ.O�@$!X�/�"��vajBT[SUB�<�Ǌ�b�$��2?���Ʌ�U)��X���ܤ-np*Lʒvv���͆��,�!=��S]������.��|�GsVzR�m��3ާq�τ� h�����K[bѩZ�n��f e���!���aB"��Û�x�6R�
��C?��S�]���GW������j�A�$�4֮���jEA��#�F�JW_Q�YyR���9߬�4,D���V�v=M�>�=��|j��ebzZ�+~! �d"pn����ꁷ�Цe���FM�v�/=a�y1QmE��Yxxq漿a`����/|ն�/�) ���%�J����w����:�޽`c� e�r��HV���h�0����4f�_��G���1����0j�{;0%&&�/#���d�x��E�C���S��I}C�����}�#YD�����u��*� V�������i�7�q���-]S���!j�"J�
%��w}P_��<���w|]n��S�q�lB�|y�6�9��$	��7
`Et�!;Z���s:�5;b�Z�:��Q�D�����ӟ���<͓�*a���c��g�������(�h�Li��V�5�w��W��C���$�Vp�C���΄�Z����bc�N��/cj���F%C�	x�|����Y���!n?�)�+w��޸���<���42	l�J�l�AQT��k��0��ܘ�.a ���% �x������M�w�=�#�~ư���k��ڪ|���ƽ[؍qJ���� �O1Lc�T3+�K�u�ؗ:�N]��cD�umC���Xԫ��=C�\A�MD��A�_qЖRD�В�"kv���G���>>��ĩ���%�ޅX���O}�Q� �� 	�i2�n},��:di"�#Vu��dĘ'e���(1����M՜WdGGK��/?�ج�C�19����C2�����m���e	^�n5�>�x�#�$��/��wi�E��0���󋘃��?yl[�dR�[Y%����$����k.ܼ���MC�$0A\;��S�L�t��ưi[)s��M���HWPP�����U�
����KQ@�܂q�� ��l{�}:�k�"��` �����g#�@�ȑ�[]�Sԫu�c�����Œ��>&��}R��'RW)��Y5���b�]�	��C���JV?����"n,��j7��=�\5$1��Dv�&�I^K���M2F��Wv_и]"�	���2SЎ|����Ew�֜���қ�g�$�Ӹ�m�(���s{��R�ECb�/3�x�J�$F���J�����uH�u��|����j���\d��A���Y�r����8Z���J������v-�_��Rh�NPѼͤX�\���ݜm���c)3���c��;���������.ڹ��>揄>�&]٪d���FIuEm|�tL���>j��b�Ng�5��yK޸Z�#f����{���4�(1:�%���8�_����=�5���I;m
��'�P�HڋkZ�v-\�u�!4""a���Uz���:��M��#��~v���J���.6�KKt �C�\�b�H?��Ks#j�(�I�Յ��RNFF����-�Ĝ�Z�q����2�߫ݨ��Wͤ;4�+�������V��~>h7��k�Ң��r�J*6�I���1�Sn��S1�������~+�.Bm��M����S�uJ��׶�N��;����#~�.n�<������~;=��<�x��������n��.��l��c�;���y��HO/Z��UK���/J��oY����i���%�w=���7��cT������{�2�bs��]��E�Έ����@��9]�?z{��@��r����N�OŮ=�9ۂ�>��^'�uB���u^�q������Ԏ+�� �.8�*�$��o�$V���8��ʯ�NO�:�+k�hR�lB�!��~5���=7���w^�
���Qu�×^�;����e`���^`{i��%3l�n���'&�(q�am�A��6k�V$ ��8 %wn;�V�̳�����}|���Z
@�G���u�����ป�_e��x��� ��Z���t��곯�W ^X�|L��P8 0�ǫ�̙8[>_���.��Lj����ȥ�d�@=οa61OH�R��_����r��kbIK�J��;�����/����w�d`o�l"B�[qg~X��Ki.�����0@��o^8<ɫu돗���$>-�g�!LRDjXvϴ+�@	o���FI	�i�y^����xnf>7����t���V�����4z��R:[����D���6X?�!���r�ʢ/�
�ƖB�P�������vY���vP�M���9�������:����h���Q;��|�OO<�sx�dm�	�Ɨ�F�_��t�\�*>��34C�H3�w/ց���o����#�A,�]v�[���#_Y8��-qb���=>��CG�QrJ���м����{���87�w'�+NBxh��2^���l�=E�bO2�'�B�)S��un�(̽e���;��;�*�yZ�}�ϥ#Ę�n��

��O�g��cc;�8��;���Z������|��u�=N�&b��{sZ���6������Iol����Q-E%%
�-f�(�	=��Rz������|���f��=rg'E%F�~/����U��k(�ۑ�����.�&��)���9��<<��W�Y� %��8́��F�<!��%�=z�����F'S�%Jp'��K/�8�KJI��$�0��d?��*���>��S��1���s:�[���A���}��/�w��DE2�*#��Z�2���ʱ��֨�^s���[������Bl�ջ2{�	���%��l�uǂ�%���n:(�tD��������C�w%�N�z��(�ꩩ�jU���`���:p���l�|�=E�~����P�U�\�)9��Y������g0�Q�LNV�q�����W]��J��?'���ݴsS������gf��� ���y��eg�s!��/8�.����꒴6m����������Ӡ<�-�.<�p�	�;����մ6%�ڶ8Rp'm<�X���u^EŨ�$a����a�G�&U�|�C�7�2�/���x�M\�U�����é�4�Rl�On�IX,;q,�zBo,[ք̵�z�?��/��u�҈��������ޠ��^ ����%�ǒ��G���$�|�'�S�l+� �Ó9h~-���sR�?@���,�l�Mx���T2L{��Rc�9�Qy��x]��WV�Uo�H���B���hhi�2*��Z�ir;�!=sGz��RJg�.�O���;�W��l�	����y��=t(>��È�3�»w�&��BB�W����/yoc\��}��r����G��b�������N���S�P�>Z��˧�46N�?i�IR�}�R�`��Fr�6�to",�8\����?��纐=3�k���y}��*$䵗����#�Ǔ'�5�d����8���W��)ݥ���ѼSJ��aGx��Ir,ED;�����I���C��7�X�����W��.Bˮ����b����T/d��rp���t�;U|\_/���� ;A��cc`��GeR.A�ov��d�y�)vH�Fiz׽DK�D����L���i�pi:�q�ϟ?�J���yOV������2�E��T(CP�7�Z���Ozj�������Q�
 ������=M��Sݝ2Yy��]���j,�Ǐ��>�>�w�{��L�^N�nk�F.9B��= ؘ���↘�|ܶ�k��F��u'�k�V�[��f�'�$m\(��`�m<�%t���B�{03�_U&�8.��h�A�� Y�ˀv81�z�<�(���}cƺ�QZ����֤���T�yӳ��J�Td���gxcdw"VXNN��ǟ��b/�?��R{��O�ёǽQ�‍���Q� 	T�T���;(r�c���� ?Y0[.T��%��1�t��e��Hz:��QC�_��ͳ���0�wZZk�I:5���o�T�XYX`�����U���߫�t��%�GMe�Wl9^�|�5���!�����Ru7m2�)�&ks���+�Q�<t�����6�(7d�A��1�����+t�ur��m
��W;�����|�{���� ����_f�wn�}�!��/(@ڨd
�k$��()aifw{X���V� �av��xh�%m���P<����`�B�l���<���>���kk��z[�M�x��{n/8N��\\j�[�p����rb`����R7o���'|]�.X�m�nШ.]�TdMN��Vo���u�O�g>��/����4e/����q�e�_�n�|�o��R����'�Z�K�͚�򌠂�	�p4�����_��,�K ��$H���e�V��k���!����	)LԾ�U?i�hC��MU�y�
4�bׅ qppTl�L��S��.��#���Q
�_Y_+t54x�+����������5h�PHa�9�9i�󺻀��`Q6��ဖ@",���_ c7j!uss�zt��h��@"bϚ��Ӏ�N�����v�$|����O��vs2����̚�fC6C�:��\x<���s���|p�ͤ��F\LDfu2���"��P�]zHW2X�(��_I6Aw���p��ap�
�v4�|MO\'u�]H��~q6)�Ŋ!ٺ�9N}�B���O���"_)�A�n�B�.�肵}715�ݽ�h&��F��,�<���� ��9Jlr��|h�I �;n��Ov��?5�d��'� ~�DAE��M�$� '������E����� q���"H�T��c����͗o^�*��Pq��[�Io7���Up6'%���')l8'�fWSCEC6񾰰��P\�4������x���yCw𥚎}(�3��1�.�����m��I��cq�	�g��D�H�o�om�3��e��#�T���M��*��B�N4��ݯb%.��[�^WU�AH� 6C���`gi��	�s�ϝm�U�c[�A�6! L;����1��+~tC�:�J�����*Pd�? �Ԅ�>ָ���1{˯��0� +�O������B+�Tw�����\YN�髁�g����C������,������:aH��!/,.j��y���b�����I/zȌ�'�۱7M�b����%5Eǹ�ǹy��Ff�[$��>'��DҒM�o��(>��o�/��Z+I�\>K�/�O)��+ȱ�$��W{ �e�\nm8ɿ���E���T(���w��,^ ����h�I�Hgam-!Q��3���e���-,?�~g�{ f`� �Ė���o�?��Z��P��~�Ȑ��aS���bHB#F�N�^�Ȱ�L�E�.����M3LA���`��L {t�"�[B��{�(�n� 
��a�"����]H/�p5\��'�mE�L�uS0��h��`�u�BT��Ŵiٲ�r���Th�1�d�c#�pk:#�&H � E\��\�(�N>0f��?� .o�كOlVÝ;}�5"_m�q���B�ؙ�~��T�a����K�z1S�������Y���y��-�l�֋>���?8��gB�n�D+�cɀ��6iИB<J���[�w*�&dX(���z�g��U��'-��>�f2�.���"������.|����0�0k`�N�	h���ð�������MOO��٢aF�6
���ű��6E��1z|�����?M�络ɀ��O[\f�`�:ۆh9�x�Q�`�g��2�!��}N�4�F:
�:��z_ZzW�콼�yh�ye������n�Y��} +x���T �.ŶhhkG�Đt�^� ���t0->�\{�D�x%��6�@-T>���ewP�����'c�?��//I2���pt*�:���3�K2��(�{pၐY��QI$�X�{��^Ө�}^�t����211�+Ӯ�7�ɝJ>x�����J�G~����C���{A$N�жz^���`gT�cW�����χ�'��(_� �*2r���,��� d�M~��_�<W�Zuf�!kG��zR��uz��5�x�&�O�p����u��ʊ�>)2T���+~��7�� �;�1�z�2Y,(��3��4-Ez�2;!��Ͼކ`�|�Y���C�v���og9��y�s�,uaf ��;�͘c�q�\�Ď��ǂ�$��H�M�Ae�Zq�s��z�꾧���p�U��SV:$@U�쪾��[��Z��ӧ�OC��L_7r������d�����|-��?��{ÿ[�KC||p9����Z#�o�\��	w��:�XV�<�O �f:�j���&�<��L�,�
n����6��K�
+�-Bm�8lϜy���nֈ�.I@NC��;F��W_�a�E_�����dN�Wqr�8��Zq��wvb���֓L�A�mVz��C�H�������#~P�ٽS��;�cY�%��v����T*��$�מ���t��O�Io9�0��{[L�����)Pʐ�q}��������T.���M�i�k������	,����48
�$7��F��&}?��g�`�$Ӈ�N(�3���F?{#	m�&�G�Q�/��w�o�~���
��Q��Er;���1�M�$iiY*K`cm-el�d�Z`�dfG&���uG�2d�,���&�P�ĸ�_��N�Y��A\��`�̘�l����x�z5z.WDDĴI����Q�h(!iPjm�_����@l,HQx��6ĩ�g) ��W@I+)nr��Nj=?=&O�����嗕͘��H��13��0N�B��Us�K0pE�����oya *� ��#�E��N�g������M��e��{&0�H 2���i�N���S�U�fl��^��;aA����ѽZ�DzY�H&��[��h�Íd
�'� .
�R���ihh�P���p|ײ��vj���=Tl �����^�_�͖
�l��wA�>PQg�2l)�rɟv�u8���O+�އ5s�h�:�D\�2,�VE�ۭ���0�V�PN�ل����X��8�&g���iK������uu%7C����XE;Jr��?{�f}յr]=&�z�
�� /0�����W}�L6��� ��q�6~	�А�[|�P�����Jtm���Y��Z|����`�:��.WU�y����V���0�Z%��Ԩ#�\�C#7�������� �v�rc�`�{>56�ӽ��O҆5_�������塚~�|)�����vL?�^��(ϟ��>�Z�I��ٳ�IU|��I,9��%B ֊ҍ�j�ćJ���o�oNM��p"4޾5ӣ9Y�Vaē��gχ9���b��OL��k[�]�uL���n-!L��'S���HK��5�=��=�# q:yT�h4rA������r'��΍��U��l���"�8���!�����9��qN�8�kh?�+���g��K�nԔ,�O���HO_m�~D�����͛-�N��_PP�?^����d3v��y{(���}q̒���ɠ�����c&��z�4$<4�����|L�󔶷��1����2c�[��E����������t��?�қ�n޴,6�G�V-�	�P�0��q�;kI�;����~�f�`���$�Q��\��߹d^��k��K�Q�pU�kkk�\:� ��A��&	1��x�`���&���O����W�Ũq�mMf�֟b�1�(��k��z0�B|���#p�6.�_�=:�i񺠔��G�������A�6⹸����X��6>K��Z�U�K��0�֊�Qgz�&6J�lU���S�L�v\,����dIX�}��=�`������t.�YǙ�� �m
��v�F^[��<�X��Ko�]8�P�Ї�1�1T2M��o|O��1�o�=�BP'j]+��y�`7�T(��T��7qtTT`���rB��^�e�[����P:Z��ckN�_$���.7v�?�^�K��� # �*�:�㕝*����n��N)�܊���֙��I@�6/��^D�:�u��4j%g``�lz�m���!|. ���;���2PV�^�^�C
���!���>�LZOa�A�;p {����ūsJ��� �#>\�Z���PEN���u�<��×�^=�5�g�	*_�M{��^�P��C �0�?�>�Gkyɹ�fM/.Ƭ���'B����2���8����c��3�wGxd��4c>���N)��߼��� ".&����,̩��F��J��<L�"s|��f���l��N���r�_�{{{{��:5[A6p23ix�e���eq�p��w���+�,�Ep'\������A{Δ���:tt�Q�H�� �:~%�Ҏ�!��@�Ѻ��	�?'��_b��IT�N��~J�l��y.����r�B� V�2����" >�ޗ W�t*+�W����z��xC3���R��k�ߚ��A��zl(�R�l��&?�:�!�=Ի�J�'|@ť���nە�'(o)���O�K'"^[�o+'��X�65�}-~�(��@��u��/�텽��L)�O�=��8Oy�ǉ�O���I5ޖ�osLĞ���ݔ���]	@�x!N��b������Yv���"=%��f��E��jI;O@��K#���8�e�;x�p�K��ï
���+q:Yt8�@P�Г!\C��k�R� ���K����p������UW�����ٙ���f�I�uG�11(�(l�0�zyy9C����]�ϟ?zN�@S?�����>ۊ~>	����RB-O���29�����xo���akz�������F��Pk�_ �4��3�f	�qǬG�J����h��1HI�0E�4�X�L.�f�p2�G��&%'�JQ���y���=�U�jط����x]Cø���əX[��	�Ҙ��qt+!A�y��)�Dɪ�1���s�;�_~��N|EJ|^
P����j3i������Y|pLp)�g@|��~
�-�<��>*���)96�Pu8Y8�u�l��A4�׺Uh�Ʋ�g
��D�r���Դ hǭ.UqO�N�?L�;��RC������)��j�Ԑ�Ⱦ���>
"9���d�<�h<�ܱ�p7�*B�jI&�Io@�;�%�:\��$)"a�'&~�fec�6��I��y >��[���p��������H�����?�������F+�;K�	1��M?����c�: �*��?s�s $))M�0_oG�y���ǏZlcTʪ�5�(�5�Z��!�~�#eg`>bW�>Cx���/ڧ��8+˽=��g>T@tgt�h�~+(@�uT����gn�t
	�r~~b��>�u�޽�k���g!���(��^>�Y(��8��t&�<��2�D3B��jI"��W�o�u�����m�f�"��
|<::Zv϶x���j_]�I7M1%�#���ę���DY���ޢ�Y�=R�������������}�+�V=�{%I��=��������J��ᣝ��8���	���t�_�hղh�BX�fpW�[���Gm�I�3ƒ�mr��Y�U��XW����W�� ����N)׬o}��f���X�~����H�K����B�h��0$��R�W��Ot�G[�b��g���؏t�9غ��PX#2���ٗ��\�&�k�J???W�Q�4�����I%�}z���ǒ����v!�Td&���(�F!Z����..|����֑���O���X(I�/i������+�SJ��r�]�?U�wr"a'6�WN��&�H���~��	���\{"���?�����_�:�Y���Җ.����h��a{�ژ��� �y�����옓���mo�䫫)� B��խ�T�όe�>�c�a��vd������ �q��נ!��엫���8�p9DҶ�=f]�6�['8��3D�*��^��=p�/�0�to�㋥|�b%��H���pQGe)P�~���= U�dC ���<񰱱!�[���0ѵ��1��7������-��;2֠�a�ЋɆ�� >��~�A��[���T��jHv��(�c�)�&��KA)�����k$~(�����>lm��6�[����p2Ӂ?������HM.�߿���Cp>�R?�� 7�[��P˚�#��>�]�X���	Ϸ�#��/x����.ӊz�����B�߽:WA�q�aPǮ�q�bwsy<ୂvZq0F~f���'5�����c�B�����I4��?�3'JG̺�[Q�A��a	��)伥n6}ju�V��"��$�kě8S�v�0�vkk�d��?V<���M [NB�Ԋ����͉��;6�v����ǍC����71"�So�ѻw�6^��:��3�I���-�@��K��H����txq�N�sՓ3�p?������r��\/o�
`@icgg7��O���V0F���@� �P4[^_?�t�77���� �4)�����Ծ�ǽ@G{���SS��'�v^��G���.t����B�[�^�@_��|��Y����`���/F�O�Cx3�欢UG�ĥe͞��̴��WaLƢapXX�X$��Q�XNت����)&��eE�é����9���M=T���΍��Iy��`��	A���k��f�i�op�&�Jo��	��F�(qܞ�l��D�8���j�C]:Y)���f8_��L�1;+�/�0vw#�d�����Q�B��ߒ�j�t�$�����tZ�n����{{�/���ǀv"""؍i���7��͑Hp�?.��PJB�j9.`�h;��0%�7* 1GJ�J��Xsb��NƉ�����_wL���1��c�|'_&BU_���,�X֤�FMk�/"/��kt�teD񊚷\��_r�\3� )_��Y�[P0\��5�����rOc�M@�2�� �+���ߖ7G����-�_b����m6�͇��,u�(�ǂV/�����UK��
xA�ݾ3�S��7/	�̬��3zB�,��7���17� ��%��h�iu����ܼ.�:�q�{mB�~/1�@
T���HZ;�E��lt*�<����ĹOJeҴ�\�
�h�!+����=E�����Y���Y��q�sų�&����}�g	ކ܎"vz���3����jfD���5�"ʺ/B����%����d�n:���NL���:
���7����+-���-*hNB�Cpm���
^ 2F~�~����Z�������M$���q�@_'K�H�(��0b�'�Ѿ��|�΢f~rf���z��K��4[�I{���ݓ�co���\�i��!�7mkT[0��@.Ƣ�3eY�N���h)���2�n�,�ǝV�w]�b���0�	�4��`�	Q�����efv6���@l�x��C�U�Eյۡ;�Q���NAZ:E@�a@@JJ:�i)�n�����S������w/?��̙a~{=ϳ����g�U4/�t��e����6X����Ѫ"_�E�KJ�Iu�t�oP�i,�K�Ͳ��#�بʨю��^���t35d��|%~F��[��Ǖ�e���Ҏ?�B\hx3�MdoO<�!ea��)otv�u��ʧ�#;M�l;�,�K����˦�r9%���p+E6� ��1	\9+�Ayt55���o߾���_;�����T�S�9,�4��]fB.���@��Lkn���Xy ��}$�gy"�L�4�pO�of����˹�y!���Bo1��'�����JJ|��!T����#����"�o�*U��l���$�e�G���Y���,�qRĐhB���W��9{�9�@����Ê���.YG�╈],5��;;;��bәb)���?~�E��>4���,����2�ߧ��>�ub��B� ��
cXD�%�E�9�%�3��3L~<c,�	�ktʖ�(��拯��&Ya�A�vO����BV.��H7j+��[�Aʼ��O�[�,��U��ͳXmW����sk���k<����'ξ:��3O`@�`�B֛	��M<����̵H.$�"�^�*���B����rXTʹ�V-���`2&<{�/���l)#�)C��k*�_{َ�g��P �mh�N�&t�S�>��mP��@�����D`hd�82&cd4�s�}���Wx�7�䐐ɦ���i�O<�BN�����
����}i�3]��O��w�NP�W��K[�E` �'�m�M�ˍ�0�}Q{�$(	����S��)O ��Y͸A����$6˧�t�z������@�yv:�$�k�f�&�&I�j���:/����������dz7{J�����������~�i���Eq�E�\�pQ�6�ĺ ���p}��ל���û����V-d��IBA�h��Y��wc�}��؃�V����$OV5�-�2�%m$hW��C�zTQ��1�/�Pl㮛A��G����m�o�	^��^�x]���&�;"�P����X5�8�wO�!� �;CCC��rk�k��TL��r��9���].�-:�j����Z/7��R$)�@���g��U��̳|n�g1��פ����s�,�|r"��wx���*�O-�*��:�c�=[gOΐ�xUPYISm�����>���/tG��U��y�,~�0W�G|�/��*�2D&7>L�c:��lw��iQԲ&+`�\K��]y�ryE��7鯬�YW��WEAc(!ad�(�y�)f��+��`��e�Y�E��P���w���Qըh��E?Ǥ�šwR�8�>��j�E��C����X���Ag�&9�Uߟ+jC�I��z���mQ�V�I}5b��9��v{�����m�����(�go�6n���G�ńk���6���r�Ƴ|��UO��bs�Ȝw�?�/��G)4��
�b,K���o�4q	������J;5Ʀ*�����@��nft$C$i�4|w���29>Nf������5G�a����v����˩�����S5�l>��a%Vr�7��W��dr��[l6��փ5k��J$Ux˚V����߻��H���k�mʂ:8�1x��V@�N��%9�?4C~7K>��f�GV��E�PG���A5$��U~HD�����rE�FUh̛mf!Qy!"�x��IϘ���Cj�Kxr�io�!IY�ɐ��F��D�G����7��<��|m̊3�&�Ѵ1j�b|&*2фpey9���5��K^��E���h�(d��9���р���º�T����c�<�o��$�(Vy�ǘ�++y�nM�^�k��pKR*�[>Y�����Qؙ��>Bx��3�M^�J�=�+��݌�둌�z�����E��R!q��Ҍ[H��i�y����z/� �B)Nc^ � 2@�a��1��=A�(��٬,n�}<�{�����j²d&&&նUm���$����W�3�:J��c!�V��,�6�EI6㻟��X�|�J�a��::� E������6 �:2j���QF�Z����~O�?�5�3�p�mC���]�T�ݔ��Ί���gqJ�����a�އ���_��������C����k��n���P���_�KE�Ҷ6	�G�Fq��3��U&�]h���X7�5�_�ݲ�)���[9��� I�L��d��
p^Y�����!eb�I���"_Q�����,�΁#��w� Lyk�n[Lݬ[y�7F�|�|3�[��P@qL��/������&=[��_?��l`��I2E��'ě*�e�@g��;��m��m���2�K���J����!Q �����kFYN2_n�(Od}��5V�����%�Tп*��^dUc��ȭ���?LR��;�'t�����>U����NV1s�b^�9��v���������Gd0�����j��"ҙ��#z�ȇc]u��s꧗X(1�$$Zlv^�zT��:Hf����~�n�q�Ph����?Un��E�IT��m~�SG�����R����W�n��wC�K��R�q����q֓�� ���Ӕ�k*�b����������A�����qׯ������U���V���v���-)���C�v��m��>��tG2��"F�{��Rbg��:��gL�[���r ](����[�uo������Sb��/�8��r2mlKqÀ�1YT/��^�pzydTT���Wiuӳrx��P��2���>�x�nM1w�b[^Q1z�G���U�~$!'�����9�ALY_{������[�*�fKT��q���M�o�&��n��bw��{�nڲPI�|�n1��3�[�u�.���o�_ܴ2?f�d~*���[t� �D��>M/1@���B	���A>��`���*���}�A!�1��x�|5dgs�Dp@�,��������,��;�}a*'{gg3F(n���9Q�z�B�Q;|��艐�Z�e��-Y��*�T�A+P����m��Q������5����߿⦶ō.c�qc� Ѫ����}#�<*�>[���0lu�4�����٪_��./�����)Oi�ٯ���6[ﱗ�i���hDm�	m*��K�%�,�d��3�,�=��o��m�}�L�D �T�;�*�1�oa��U�����^�hZ)�� ��9�@�����-s��o��2_#q��y�1�����$�4y����{�b��0��Z�7n�x��4���<kr�v���xG�b7���"�B�/�L@>+���#���GN<�D�*Z�)�W�h��?j�8�c�233)�N��F�$�	xZ�AM3}PaH����>�b�����&I��s^);�����.輄�=�U0��y�,�ɪ� o�立��a)�Ksˌג#+uDŗC����� 6�?DZ�m�29%%��^�}�7��^�^e���t�۪YNQʒzz,����U�d�vYC.��RA6����b���  l]�	`��APdh��]�K k'����������i�y����@�sTw��%s���Y�*Ǯ�����I���f����]'@��j���߱u�M���*<��X� �!á�J���Z��HL��Ynt�(�#v
������H�f�LNM]��;�^\��{J�X����w
���}���{���cғ>wt ��Ϗ���=-����1,Z������������7�j_Mܐ?��/<��SZ��,����I��=
����7Ui�@�X��`�U9'_ �{�=yYyH�CU�8$A��76��N��4�9A}�Q�"�q���s 9̙�;�%�OwP��xz���o��]�N���Wa���A<�q����-")s�����v��g��KxO�@�V��f�B�.���Q�s#��:9���.����\�S�Aƨr����g%�������4ȵ%"����7���"3�?j����-�M���wY���y�?�IA�ʕ���苾ڇ��wkg��{+�{��I���~xs�^���~�)�e�;U;;8��:;:�V[�>z��t�<�����+������,�Xm�)GTא�����ӌ׋�qQ|��`fy!�<KA�{���@ӱ�4��"`�7\T�.$�z�T��o��|��SQ1�2�f�N����iR�_�ψ�-��͋>���H�����~0vU�QHD����-,�h� �&�<�+r�V��c.���Px�O)?}�i��*d �qk��-�p�a�V	("s�{J��'�x���kB<�:��@�5t���5��f�����<�?M��\�D!�v|��� ��a�sވ�\�/�ݑ���S4"q�P	)�j�S�N4r��0�����>bu1����~	���GA?� �sD�W}��<~���TA��z��x~�aE������� ��W���mm�$*���/��S��ކ��
 �錏��`4<�&pf�[[;�����ގ9'~�z����pm0n���W�LQ������"�61�W)/k��Բ��:��9`1,��t�D{�U*MRP�C!�k2ﲛ+��N̩q~rV���q��%�(Ѵ�d��=wtw�jrA�c�Ru��) *u�pwFS_�9avt�>��dn�?k%�������]���y�XM_m��Տ&����ϳ�WL�e:3�Y��S�ٖ���A�,t���[D��s���Kq�"���Sn�5rG��9w�ƒ��-%����K(9.Q#�O�.��D罭W��6ӕ؃L���hUV��o�n�X��$3B[�]*��=�Bܪ+mYZ�_�6�b<c�ŁRAQѪ���9��M�"����@w�v�Y&p24Z��M����!���;�bG�Ż
N��W��o��e�b�������3�MM��
3O�G�%i�K������.����z}f�r�U��0Ta_ ��U��ؓf-�Gl�c�'����l\��68���?���%v3V�l(%a�ڂyc{\NE�Ԓ��^�lp�	�Yw��f�Y���ً�l�e ����Wr60�F�i��I��M������Io�K��v`������M�`v���̇���>����_��f$;�p�T�P�1�\���jlg0q�6k��X���&�9���$X��G���Q�KEl~+0�]6�)b���j 7����hKJK���?j��z��RY�*��az�8cpgzH��޶�����Ȅ�آ���Q��*̎���I����AL	{���+>�z�}���r|���ޯ�	#7a����WĿi� ��DuD�!`�j}�B�RQ�?.U�d�@����LlΓi>��⚡�Ƃ�������y7��'�*�F� ���o��%q��? Y�o�����&5N�^]YY�z���+�:$#���,�ϸ��h����د�zߩ�M�2
�v?��+��i˼���F=	
�_}2�g�y�d�������i{�g���\���D�����;�Vػ��k�%e���on4��\)���m����Z������h��6��P)k=M� ��������Dc~QQl��"tK�̯�x���rE��>NW&oФ��2�A�Z&s"�VG�w0� ��� 8pR�AwP՞(&�ӿ��_ۤ@ÁmY��N��2::����s����5L���\u����2��QS?9��˽·S���v{?��[nv��Xgy��A��=��`d,��}$5t���jc���tt3�c���Te(p��)O+He�X�B̗�]���d0�o���a���B`1p���[&��
��V���a��R��k/UU�Z��ᤌ;�X{��e8{�1��{���DE~4�VMM�$������TyM9j�=n��ݥ�ߢX�}��\��_R�sh�ْ= 3�
���9f	��;(��Zm+q�a�m7r��ˮEp�X^\�7y�Do��5��Kuˇ���^B66�Q'��xo�}�#�͟^Cj�!��=����J?�E�o���]ۀ�#���F�I�&a��\$ع�i%��WC3������RI�5]H�e�`Q����z����kb�K=/}}y6xw�h���WSl½�,�����I��lllA���E�(>����yZ�Q~jj�1�w���,H5��f=tuj�{�v7k��h�&TH�l��'����:<×��?���y�ȯ��;�*��Y-)!
�������ТD�a�n���(0$$)�W[�T�>���=��̹�8/M=�e��8�uK�P"N{ �74~�_E2�^��l�>��!4j��|ĲR��B��z[�&��2ss�*a�K������ � ��Ms>��qok˶�E%���U�#����w�]�%��OγWVo��Rw��$�?s;�U��!���sk�����yVE*�I�����..��?
u��0U��o����2��,�����& ���uR��&ft��ԭ�����:D�	�6"d_f!Ý���ܼ�}ie2<�QgV)=���3�)$m�����G�:���&��R��C�[o|�ī�y#�SPrbp�C�����	O�R�CܺKtJ���3�3��5�����U[�4�Gؖ��(�$.h#.Ƌ̖&v�5���s:�$L�≊�N�?{�D��͹/��qy��E�����ތH'��6Ӕ�%����8�	-T����$|�Dܺ��,�����,��" e����SeU���Ln�uә���O��imjV�Ԟ8���v&{�s��x����%��;�J����L�3�����P�x�~��/C���B�&�};����C�N��US�#~���@���S����ߪ�n>�suR�gV��W��a�9E����i�i� �ҪO_噿Y�x]
�7��g �x�u]a���}�z���egwMZZ׎�"��ԏjT��s�s\�>�++t�FFV��c2��;�Z�^:����8c*�,p��S�6h��PZф�V8+q��u�j��D�i���R1��� ;v�%�c�j�����Ԧ�ȯ�T�+��.��!��[�e��ᮽ�W���An^�:����<�-fv��\�	ڗ?1�{zx8 �<�tF�w�U*V�W���h������w��X�"$��s��vٝ+n���g��jy�ʕD��FY�ZQ՞�!kt���w(6azhh�e%��
NZ�=��|AQcͣs������hF0wɐ�#	�A
�q�"�W��@Lp��*%�J��0))il֗�:��T�GjOOS��YI���y��#t��H��I�49��Oߡ{���5X�8C)��f���GR�L�w0q�E�����h���\4q�������`jj$-�/r�rT&S���u��5��A���a��x��4q�ɠ���hn��G��;�|	���7����aJ�s�����'�ݷ�@�6E�S1s�Xbm��/Y����7::��$��������,j0֜�yxP^^��n"�v@�(��wݣ$1$F�V�u�_痮6Sl��_b-n�����!/^J����0Qd�PY��_��]|�]���b
�W5�A��'I�wy��R��J�s��O7U�pcJ��q>�ӿn�B�f�I6���Q�5���\K���%�Q��Q�]��|��F�F�� ��yQ5�Mc �o��gb�����'��qk�ed�sENUY pxZ�a$���G>Q`��}ծZ�"�Ч� Xߥ��P5���q�'�p\@�k���)N���w��Q:=tx��ʶ�w�W._�Xyx��
�C�^�A�HUg?�s�$��"�Ξi�nb��KQ�]�d��"r�-��]�(9!��?'���4%q~oNĚ? ��j+��^\6Ɓ $�"S�5,b�o�r	d��i�x�H&�0��t���0�b��2Gȅ�C��%�7H��`F��6��|���}�ԟHN���ST����L9G`��G�p3X)����j�h�f��n_-((�-���0�?}�e�"�����_��x���W��ͦ蝍��n���lBi�{��qZ�݊gk���i���%��������.���33~z��6y�b�EH����=i(���c~	���t� ��i�%	�Bf��b�[�|�:���݇��t��&7���XT��[��\���(��B�ce]���J+ ƪ�N����S��2�^4�q/�޳���ظ�z���Y�a;Z��'oY�f���퉉��_���~��N��Dǖ�+��g�Ǚ���P��<R{�&v,����C�%KR�l��K�Y�a��tВei�T�����[�����wR&����!J�l+����
X��Q�*�����s�S�c����#`yy�Oi`L���R�
M����V�h�H��Ev�̢�X��!�����m��s��VkuF��	�=c|�-bu4�>�*4y�&QM��DH�>+R[����^KL"^@�Ҏ�_&���U:��G=���]�
�h"����}�O��,��q���~O��Y?4#�9�2L�f?�E���S}�T�	�é~���-���p�1�]����7�"OY�2�᮳ �dZ-
��U�� )4r�ve��!�Ѱ�?	&*/t���8�e�Z<���<�A굱�fNժ�����c��,�|���N�Y>*�-�G&Ӫ�U�y�E��W$g��0& nq�E<��e�ϐط׃�D^�K�T��k=������Y���@�r�A*�^��� �����EJ��;�Å�͊���e��}�_:!�w%�]�gr��.�l
����~T 
�����ی�H��V������'D�ǒ8�V2��!�Y��F0��bm�9��1d���Ox��3-���t�x�U�W](��>H{��*��,}�"C*S�;���.�{y�aܜ����k/H*�|���r��@�KW�9IZ�HV>�"Ǿ������TA���c�#{ۚ�A)�Y��߾Yg�B���uwU;d��M�c��[�h�*�t;�;�M�`�p���S� Y_�!pJ�@��������=*�z���;�� ����q?��nH6U�Gxnn�2�ά���
K�.,��[�T�h�z\�P̻�7��E��k
����s�H��ي1���Z�&%6~��G����x;���[��r�fw��c�ج!!tu91f��JO9��H_?�Z�-Y��|/��[��F,��1]��F.��	���P���!@���I�����n�����ÿ�b����>_���8Yɱ���u�e�]t�l�����f��9Ӳ�"�����P���p�cr����|��Qq�5r�l��{�ƞ���!��+�`�b��6���a	<ß���mf0��r�<�����Ra�t�H�8N����aF(s� }J%�Ye�����60(ׁf������cУJ\��PH��̋$��T妚����k�A�t|.��Q�h���ꕀ��pl��FO���U�f���3�4�����	0�Ҥ �>�B��$9MOG��ϟ��ҧL	Or�9��le���Y�#����3I>9�՚8�	;�����R��3G�u��Z����s��m��aɑ�	F���T���Z o�W���n��}V� ߹o#�J\�j"mk��6�%G���bG�w��J�EFXb��͛v�[@�cng߰ͲE�k	��[v�>��g�}'>�����n�O;vv�|5Q���a�$��Ɠ���RQc4�j�蒱8V��ҀQ�bj�$����4F��5ɹ���Ꞻ�)���/??#���ӧ8N�m1������~.m+��{'�O��8�a�u���M1�N����BSR�=�}�Z~G��-�nӒǓՌ3�;���tP����:��8i��#��uu�,�5�f�3r�Y �Eb7;������B�!�}��N谏Mx6�p�(-$���z�If�G��|�44D�I�@�82�px��m1$�H�Ơ׊�U��3tJ���A�Q�xbW����S6U��8ΎvZ'���o2�������L썋pth(ڬ�@7rd�Px��X����y�J�{�~���3S�:��Z���F[��O59<�;�5���?g[t��o��$S[�r��3#�9��t�>>>��W��zb��J^Sβ0�f�I�$�6�i�:���o�~�Jb��A��~!mg_ ��a�^%M�QuM��F�l	��9��R�.^�V��q+�^��:1�Y����`�z3&.�Mf��Ɨ�����^^���h��R�kܗ�gR,$������P�iƊZuՂ���`��!�
�.���z� �� ���{k�s���^���iD�k�\n�#�������h����{��
�> h���!�<��U4s����2����A7���9�}>_���
x����%����eޓ�:�v/��^D�a.�VUU���O}�0����_�Z��l��U��󋋘��?V��Fv��T��{?N�Z�`�L�<��FO�46O��·�PaT��io�=>>��T$ ������h��\?/Y;�k{q��F>��1��9=��P�eӟ�\B�cY��l�T�h=�]�L�6��ԇ����/W:�8��҇|z�\`���j����yVm��mN�G��Y�ܳ��# (=gEzK��z��z����M��9zV\�>�D�
3 ���N�%���%ϦS�Ģ�'���B�ES�8�ܬz���uu:0���G��������>��I,�/���ާ�'Q��U �jaa�J?�Eݞe2�O0ߡ	�ڗY��Ɵ�,��c�(��#%�xA���+2ss���`�&�c��P�h�(^��6$������������^)>���_���oJ�P��U�a��ˡu,��VԪ�Ǫ+l��9�V��BM��--�0ahh�r�&�o�g;ɋ;�H�~b��ΐH�~*�7/�]zf���gIp
e}����@�L�|���.�)\|�#W�o1>I ��,T��]\Dұ���0����C���v��/y���vUǴ�l�j�~��L��"ɒg�7�0���ec�;�v�+�2��F+F��G�o�m4�]� ���7�����|8ݠll�hى\%&�%�f{�+E��7��Q�N�����dݷ�z�R���2�-�A�
�T�S�(�ϟ��7u�EmY$��]>_Q�t�%Q_q%+/�⮛lu���ڀ0��%�mpe8�C�����k�E�3U޴�|������m����D��A�Pi����Q�'�������ۤj�\�����<�����
"��$̄n�(�fZ�q��2�6�S��L·�.��5`���BjZ���k �jl���o'|4`$y�� NOV��7%1��!�O��~c3℞a.� �
��)�Sⴽ���M��ܷVa�����;kt̘�p����7~����)�/�k���QK��S|%nh��dEr�����ڝ�@���cI2슸���`�FW���k�ܙ�W�>�5�w�x�9�����!�h�s�=�A��~�1w���&��)2r���~��E�=	�(y����uɐ�%*�ʊ|�XI��,�ǧ��=D˯<|�tA�������;ۼPלge�Y�ֶ��P�_�d�}��G����Rµ����[V(�&{r��U5Eؓ��o�8�.f�=,ə�}f�����	�^������i�U�+���A}"_��ns�
K鷬���N9�dQ���層�����wF�����a����U��15�<�mX��l_#t�6�{ϰg�Q!T�e�N[婶K;b�'##����٩�CT0������KnV�{B޼�L�ѐ:��r �ֿ������ݰ��H%�@���8�d�fZ�
P��+Ziܗt�� ��1Y��LG��� ��whoԕs�-}b��%��TN"W�j?nH�	�]��i�SE��~�H��ϥ�����fO�!9��q��x�0�ŗ�+�������>�U������H�ܡ5����cP
��q���lw������2ӆ�B1t�򦥥�m�������S�H)B�p����/0�}�W��	K�&̆;p����& ��a�����}��x-�����
�6��3�^
B��ė���ո0���� ���F�?���@����_iQ�M9]���T＜Bݭ�V(=�˖���4|j�-t���VS��p8��w�a߃��g�M #z^L=���aq,��l+���dw���;m;T����,������;.����a��ϑt{�fA5]_,��n�a�V=�*=�C� ��k�Z	H��Fԓ�(�~��LB߳��\N���
ߪ�~�]�|~�z������W�=Πߑ��e�]�M�~���S;[�����r����$P~�@��f#�*�s:�r0p���Dţ�3�����ʄ*�^��'[�D��N�=�WX�1_�,�y��v42�b���Ț'�Jv��7��8��/���jEV��qO����xL2.444��u������i�M�������Ɏ$��iXt�_�b�H��D..�k#�"p��&�@�F���ݼ���pM��K�����@���c�O��ԧ;�I&8����d
051��P��(�^�Lg˧_�d���1��2�yR�D2B�^'O]�ŗ�/E���GA\{�]g�>~�Yq�Y���f�|�u%���K?�tO��Ǝ������M��~������]Yht����j�v�o�ib3��!I9Py���5��W3��� J�,�:�S�E�U�,�n\K1�ӭ���=���X� m�:}�Iv�W)�]���#�@�E����ox�&����F33��&''u��K�I�+��t\�e47"Ky�˓+Y���j^EB�S���5ٓ���9@lW](��<������%j����Z���q߳���u��Ũ�ҰS�3ޏA�-����;�!��5�k�q%ǟ%���O&z.M"�.}���'�
$Z �A
��1z.��{�Ά� ��*�,Z�@� ��@G�ߧ��aYD�73�͓�)�����˝�.Yww~��nZۨ'_�[�
�j�62YL��CV�%��
��FG���źo����1�--}
�e���!O����r��E��eG���}4�z��b��zgډ_�ɑ�'��T�2H��{^|||��ٓ#_F�R��]p���/�X���#�x�x@�~卮�&3!�Ͷf!)}O{b�Wm7(✇��SR2;�<P���J|Еb�Tr�/� C�QOՇb�N�w�!�<�?� �h��^�^�ġ�sMmcK����(yh�E~��X��*3����b+̉��	�k?��P����N��P��'�'I={F���0��8��!�%F��3�跀�'�w��tٓى,D[\��[�~�ߐ��O)��*�!�h�b9>��sK��V�������y��`�y���k���8������Q�<%�)Wo[N��k�z�����=�[,�В�,,���'��,�\�m>�kO��]WHP0L�������Ϟ;��R�|����&֜?��BE[�,|��PVT�z-fx������p4d��IJ-~�#BӼ�q�n��M��i@�U�]��9����ؐ�����k������sS��������h��m�cc?��j�#����@z��j_Dސ��I�Ƅ�K��	�%Be�\�7} �,4�"FY�X[ki�ag����Xx��-]ʻ[pr/z����94����Ԛ�s�/��L��&3_����T�5_wc�n K�p�N�n���`!7��m��|������mɝp�s�����ߕĔ� I[�89�$R��
1M��ם�gR	��`�a���9ŭ)�j���|��weɋ8�-v�3_���z3��X��NNj@Bۦ���*��`��k�����
��:!E��?�@��\y��v��-�	X�-�/^O�ۿS+��=w����:*4���^&�h�St*'���ziAO��2Se����B�U!'�^g�W<+�%�.�]1��<̃}Y��#/�m0�@�U
�ȭ��q�C�2�w-0#į�ڟw���H�,�k��*�nn�n��U�n�Yf V�'P���'���AA�ԩ܂4���/p
{��\۳�����m�+ZaGd����b����F�-��"����j�'L!R�/���m��g���;ԟ��mj�O^���\b)���ﯢossCx	'O@�d%�jpߊ�,�7��5)�_{�ް�}BGw���B�(�>����{����{@E������0p���]p0v��m��s�
=���e����H ���<&�g�d0�|��%��|d���e1���ON2+���o���l��g�8ȣvŚu�17�tll|Vjq���TUUA�X��#����D}Y�`�t+K�g2�s߿�t=�2��`�������)����:b�	LT�M7D-�}��@�������AR�u��KNn��4��?�%�+��/�y"�P�Bg\�v(�7C,zЙn�dD?{�]W�R��,�PU@H�N(�cE榮 Ӊǧ��`��9-һ���2Ymk^q1Ve�Y��q�D6����rA%ٌ�Q�Pש�����,��B��5��9���^���L.��G��B���d&_����C��J�xye���S�=?����9���|N(�ǘ4��J_͋���X��j��}����w �N�����d�JFFֆ�\k�������!S�I݈���C8�76��ԣYP��`�K���:���q��#V�w��k??c���)O�LZ�ﯩ���ۗ�j�����*\�����"�e�:���a��M��|a��a��t�����2�J�v�>������Q�錰�$^�'�=@L�UV �6�Q|J
٤�0U����bS����^k��ͷ&>��P�������aIN�L934�o>�®/�:3�ɀ���J��y���+�n�hI���Y�2X�����\=��RoZ�i��"=vʫ>���g�GD3��o=:��T�|ܳ_F�q��ez5��Y�@�O�G�����B=�[���X��1��q���]�,#҅"�р�ג��6�F*���ŭYߦ���	
�@$�Q��lؓ�#�ϟ�||�X�?~KG��,\`�j^�2����>��e�c���f�P(�;�E��(�}M��h��¥o�Յ�jY�Y`*��i�<�����A��A��Xv.R�j`"�9�-`JR2n-�{�^�3L����`�\c��)�<$ ���3���n��.���5
��甙�r���%�S�4�cm:a�ԈT�iX�Ȍ/�}�f�������Ĭd$.kA ��$����o���#�n��ō0_�����3j�E{v,F�o�#���ёT��_h�>>L�6���ϊ��|v�}��<�,���{���(?�M�s}<Wv���l`��0!��v��;S\XJW�7�O�&A�>����RT+<A�
�ks0��1~1ɿO&��NV�@kU����^�a�Vl*���I@@` ���Q }y����L__��jxʾ�!��ɔ�WLտr�P�F�1�f��_1��mmlm~H>�E7�@�����$N���U�R�z����_Ljx]�����n���,�]��ʌ�J����쏙�u�Aj�*}x:"ڪu�!/��f�E@ xdh����:2��d� N��!k)����(��������}ˀ�;�w�����M���iy�c]��u_��	�ps��f���w�X���[����%�v��S��ұuT����2$�@�#0]ȹ)㣄|�&b������_���=�~G��0��+!q����{o��q�sӏ$��^�R�?J������,e�Q�T&�6+���l8��`��8l7�:W�l�ً������QM��s�@�uٺ�@}�x~umF�g}�j]P؇	n8ccbV;�v��՝�y�n_��]�Jd+�_�������KC�<,n�[߷9D��X!�B�����NK�*׀Er�y�a���ק j!q�RW�m��-O� ���ei�[�QeM"��?�U\{�����8{g������F3��@	<~<+�����?��"���ׯ�q���4d>��dRZoMܖ���t�������+_�ȿ��J���i�'v��|��<��	�E��6#`�W������D��P�e?�#�Q�f{
���w6K׏�/S/=�~��~3_�*0bM�&2k���ޞ߃�V/��"����`J�ӡX�(cN2_5&C�.�`�<<N@n*���L�=�
Č�1p�h�E�h^ݼ7Z0t*	?os�Ng��G��<��4�����I�cX�����T���3Ѽ����5@�W�"�l�Գ���ɢfϖ�xq9�ӖŰ��N�l-kO'_ ż�k�[��"U�m4��N�X��u�a������| ��(��׾�8յX�aB�G?0�$/�>�涷�&+���C���dD�T���L��c�{���@H�;]R�@��^qj�=4U:�h5�_�������g�4됅v.J������� ��o��o��#a���.��(�����b���#wgj��O�wV�⤜S��e2K[�]�`�7��a�1sZe��1g�۹&���{�)f�N|�jy����"��G^}���b3����&���C�^��lDa8k��**W�|��ު�@�`�&҉83T�k�e�,B��k=ֆFF������6F�����Ͽ��T�Ԁ���A=Y��6���o��@
��C���Gñ+·pN��8ʔ��<�_0i{w��*��㞾�!u��/�>{)���1�T��u��rrU��DU�t��wr~Θ�f����x&�{g��C�O�b�
2@?�J�0N�A�X�^��s��O�]����S��.g����*��������h��B�Y�vv�O_T��;�i������B����0R�I[�o�#C3���0�ɚ�l��n^��5�G8����8콜N���?�P��,�}�������ڸq��L�3ȻW�d�x�)�h犄���#�IDC͠�k���r��jkO� �fEt��6HU��x�M�����exl��3Д��R�@�[�a��l�-Fƌ�q��6�kHZ�s�$����l2+jXntW��n�g�da�c���	]���X��5Ԝ�NE9��s�v���6�o�(�f�x� )�O2--q��ޞӲSS����ɗd9w��7#���UK:���*��7���$����/7a�:d�Q#=u���\o�𴇦<(�щ��,OO��<�=%ȯP�;����:.ʠk�niIi�AB������{�ni	A@��K$V��������y���ta���9W̜33͹�W#֞9N[&����*E��@�8�X��Z��7%j�(+������a��ʸd`n	�̓(����nB��`|>��N��u+q{�3UR4�Õ��%�9�J�x����%!�^<�:lK�?x���(����!�� f�r��:,����o�mn��f�g���D��_�A#bQD��N7���i�y��������x�:�����b%i dzr2Pq�^c�Zf�?����Y���7|�ݩ�/����
�mk�S�þ��}!Q�*of�e�?�P@��~C�E�tۡu��E6�;	�k!j���8�ߧ���Q�g[|��!(�ZA�������s�,�w6��& ������Q����iBޗ?���~<˼��Aq� EV}0�
.�[��<���y$y��Ǿ:�#0(���� ����x�L �l~,4���?�B�bp�N���8@1���-u���5C��/0z^$O�T^�nL�o����n���E(E�����!��	���S/����}l��H���ն�☒�Η�R�N�a�WK�܁���?7�}������#����d&S�)?�,^;�0��#iC��}Y��uI/�efrF���N�NK�R7Y�l����Y^w��@����CQDm� K�6=(>[[�V��y�nӒ�h+�_�8��Ugh$�;��r � ����]9���n�����'[�_��|��U�9z1�V.�$r8p1@z��{���f�E�R��+����;�����\��lV���FxQvpH���P�V(�X��B*cGk!JW:NOU�
-�����n��?���l��Zv�R�E��%:N� �G�>�[�N������O222��b�q����
�X��ܪ�R�?��Y�
�O�ex�Q���^�3Í��\��텼��oSi�ؘ3+��)#f|�\���ڇ��,3����ղ�QbT#��@������N����AV\ύ�����Qdvf`�7�33�`7w�f�~��`���"ٳ#zE�o#�Edp��n����i师.՛�,��yu���0w��/1EhH�'�MU{B�(�<#>=w��N=����^}w	Xj��)�m�!�f�7g��~�u3�U���gY"}���U !�Tmo�>�^�{�G"ܔ鹲�p���	Q�7��I8�R�G��\��NͿ����\������"��ÿjh�ѕ��rH���vԶN!,v��������A��
��9)���.$��@h3G?AO�����2̗9[)S��c;�{!���B0,D��$���w��-�<p���`��`?�`�Mr� ҴA(G�[G�f��i��Q�vE�N��&ť�ϝSߟ{�JU6�I<� ,�Q{ɢ�,��!"̍lZX�T���ݵ�j$nVD��dLT��10e�뢐ب�pī0��_��ȳ�4���fs��&�قT��dҊ��w �G���8Hf��:�A��7sK{�F �	Ʒ�WF��M\K�Qw)A�[qB&:���v�_ld�/��Ǝ'�x�� ���u����C^ڶ(-�� rW7�r;��S��G;�#�B����DDD]��J5WaL1�cT6Z���(=M祒�e���O�cwW��P��?���q����?/�����-�����V/�fcSȊl�逩����S>�����S0�V�� +���`�q#h��o���/06��خ~�l��4H":�@x�T��K�Ѐ����ג�f� ����f�0M�}	�,nٟ�PЏ��(�����X��o�p7ѧ�P����l8�a�x1�J,���v��	�=X��Ђv��L��)����p�KFFb|�F�$���a�j�;��I�9�!qC�\۸�Qs�	[]���3�u��s�Wy��3�|���2�����s�TO�U5)���,��E��<K� �Aؕ?�&���Bq���.
pP��� ���܌>>��B�M�AE�=]�����5�
�vFʘ'ˌ��oO���¢�<�WH�VOFU��D
�
��j��\�u�Ӻ����yk1vRABj�����m��:i��2�`��j���dz_�ت��ֹ����3���ߦ|��:�r��Zcqq�)�n���?!V��M���{J(}ӭ4e�5��m�Jղ+&�,�0`H���/者<7��Z�}�0)Qۋ=���+Uc�����n>�#�6�_�tD<ś3S��#z��2�p�c��·���ד ��I9g���+���a�J�Ah���D3�7_RJ�lgJރ�S7mo�EUII�_q��
���Օ3#c@�Z��]�/b+/<�4i�X̢XSo��h�k�'�*7�Dȣ2�oZ~g���:���&��1�x��j���b���h��%�g� �5��K~[�K�G?��_KI�۬��UQ�^M�fO����f6S�&�]$��C3a�Y��{榛�}2�Eo�M0��=�a�[R:� ��dT/������l���;_?�"-�jN2��������E*l�CJF&�m-���K�Q�0ѫ�3�æ��#�TUUS��e�,~�9������x��#N���봨D/켅�|웜������&6܈��
�ML�G���>�і����T�>�Fq�z؛*ӂ�΅�K�#c}���TaOT���m��K57��$���̛���t���&��y���܁9䚨��ihW�̢���b��~����!s���I�Pr�uj���<�U��g�V�#�D��w�T��=�Vu�GC =P��pbLY3��h��,S���#lT{J,�X��%�����Ma҄�-ɖ�Ӧ+�+3��|�$՟����M�B�Exi��}4*#���d`�ZUr񦣤bs����馘�� ����K^n�����-ڈ�A �S�.���I2�3(�����loۯ��g}�.���NP׿�Y�"�����84�w�o0�"/�j���$���&���-$ue��67=���0���Wg6���e��|p�5�a�p_>f&�Wh�R,UM�X�f�cM'Erp��F��am�Г��A�XiqsíF���Ja<T��p|�T��fC]�~wU?aͮO��l����z�*���%j��hF�>~����ى,q���+��Ϗ��a�gXCf3�!�/��e~9�Dr��ˊ�D���J���M.�p�V�������α��(���3�1I�3�h�1�K]CC��3�ml��뛚���������*1C�T��s�q=�r��Ih�c� ivf����~�B����gl^�]pj*���Č��ۼ?Z�T�W��1�׽|��5��W]_Wq��������Ō����X �:<��˛*a�ozL��L�_2��fL�+ھ�Vv3f �yByjj�2+�錴:FΚ��t���|�}TXs���kǤۨ��<pf�[[0i#�/�P�8����|��o�\����Km919򨃮����-]���� 0�i<	��!yV���E-�/�H �����`�M��
�1��r��C�:q�mV����2�4QO�tś�v�\o��L���]肂.
�Iw��*�	K��S�ݒ�\jR������4��c�mK��K��>����$tY\z�jl��uX/�-HW��u���z(eнѾ�${�� z4+���II�@O�yt�GCdf�f�����º'�V��.$��w1]p��k��h/!���.C7�m��J�FO��^���G2�	�	�#�x����"�M����%+#�'���r���e�=7Vu�2B�4+�y���|�F-�X�E�"��B��d6E-�y�����u��F[�8 h{��7�~�J���E�P��sr�(��"�X6����bw��= ��F.�`���	/��[9���J����[tt�-������}w��B���li����,�ͥ�E��=��5�>Y�nM�X6��C��\B�D�udL�&�D�)F2_�-+d�����-��	<`Nm�ǲ���%8��2�;vgׯ./�g��xy��-)�d��q�{E�A��}-|b5y[�����CG��pi�rh�T�$96$N�@1�ⷚt8G�w㣢e3mWo2�+�/I0ȣʲ��̳=qmmm�k��+��S����z�	!��i\Ɨ��O�4�)"��&����-&
=�8�����(�5�)�o�X�b.T:��i��(C@��ՙ���u�E�Em�4�m���a��T�:<�܊��4�b���b�JJ:q&�E�F"	b�v�+U���J7o�:�|Ӓf��뭡�̈́���B�mY�[.�ށR[��'�Ч+ ��ɠ�Aɵ�~�\ta��H'7#��l*�Ŗ��
�� ���ύ�O~��Jc��vT.]&����M������o�FO�D�e��ߛ6��=�u�[~��=(	���-ӡ^�vm*Y��\ڟ\�i5�����'S��܆aooo,~�C>@ �}�øV�I:]y�f�1'�RrہֳO�p/d5+T���s��r����c��L��k��|o�I2��A���4wr����f��7?�ё���	�O������̜�֓?��;�M\g��a���ō�WhGL�(��I�Z�9�x��[~�vE2����O	U�B�� '��ٶ�ːP�֘�Y�?7y��r�(�ڻǬZQ"/\���?�h�Uk%�ufdf���A���A�ma��j���Aј�8]��z����~wz�O�M�!�w��o�	���"**(�&��:&��%7wp���l�����440"u�������0C��*.��B���ƥ��D�<lh�I��;U���ҋ�Zo/o��A@�Z	��G/�Y�ɞ����-���]��-7�U4g��b����/�5c��:�D�Q?)۸���oB��c�K�����$����	æ����D} &�x���6��3��v��_lҁu9H���B})����]1��©au��}:C��&�&�e��$ųM�'&'��L�ց��V�b��oqA�f;���0S�t,s������韛���VC�����:@����7�|��|�u�/Q`$�X��R.t��b�w�D�T�V��+E�*[�G/̚ϣ 9����sٙ������6E��`yl�u��S��}��D�_dE2??<���<:0Ak�#�����1_:GA:^��d�������N}s�ˋ'�ty5����0cb��`��Ľ�:N2Z</�zrv��E��㱔�	����Q�v�y��ďV��Ź�c�R�pq�\t��v�eMK"Xa�|�� lެ7��d%��wT#�CrֲG1b�8�`�����-�ջ�1�5Ir3�������f�SՅ�$�7y�	dC��f�Z/���m=n)�L���;���r�>v�����f*�g>��C�R�W*7��H`+��n��b�
��b�E����\w�����i]8���+L�i(4�T,<6�T��8,vrwg��y�)��qP��y��GG�]\�ĩ��o�./��D΅O �������St�y_����7���-$1[��H�-@]e�c�ߏ�^L2?���!7:\�S�h�Cj�mx�3Ĩf���q-��R;�f͙*�:UB�}[��gm��e�4t+�WX^��	��>0˩c��fJ-F��my�l�!M�脬22u<�z��3y0���?111�U݂%����E����/b�s�6�(h�ȼ�҇�r��p-z�+?DJR���`�0��P���Pc-��zjVf;ǹ�}�ޤ����W���i��ߨ��up0�(�[�K���dJ�Ƒ�*���)�]��D��툹���͘f3hD��̆���P�p�Z�x^���Y'!
B���n-Q���4B@��^�NՅה��"_~�������F=�������8�M���Z
񯕕�	�zz}�~��<�l��q1KR�J���z�;�Z b�C��:Uc]c���)B�:�Q[�i@<�����Qsf��꘻��;w�vn4|�M��Lu�<��3�^v�go��B2C<L���`�;���c��Pj'�8�����%��S�-������D�t��6�������֏W@B���s)()}������Z��5�C��7�^d-����'�L��Qe�9E��d�P����N��ݽ��d8a��q=�강͏�:p�ϩ=n��B�x�������-I�4����x)f}0�@�U��oTC��y�r0;���x&2��.�Y����f|��g��S�χ�#�m�ޠ֗�r����iKE>ߓw�������آH��s����c�ڪ������N�a����e6����9�����G�Un-��(1"�p��snS�x;w�2�U8�6�}��޻�f����vo�f�y�Z0ڥ�Ѷe*j���f��Խ3�B_�����{<=\Ac�J�p�"v�Ј`C�Hu��$�+>���fs6�N��.��m>sپO�w�[JI�'������!1qW:�MKh����BU��ƣ���O�^,�'s��_?V"���X��6K��M��G��l�I�!1 >M�����p�pꏹ9�ǋ��9�%"Y���c�_���d�}[۷j�VaL�t��L�.cm�Z�Z��Q������]h����_%��^�����ۤ�QUU�S�� $������q�ۻ;��A@��}%�A1�iA�<rX�oqJ)�]�V*Y�L�ܷ�_ǁ�W��+v�_)1!���F�K*�?5-��"�[,*�K���FG��Q�ՠ��2����E�ϒ������܅W&����ִ���m\������ￆ��5��Z�"���Ͱt^j�_h������a����6��ʣ�O��JK��,G��Xg,08z�G���:RU?d�	n=�L�Z���!S|��ZC��!�ښ�w��
����D��֨��κ�Yڋ��ۓص�Eiq�G��X��pv��I*}ܽM�Z�rh�WFU�f(N�\r��:�c���8ߜ�>�X�g^� ��_����h)r��f��i �i�yt}��l2�ܪ�̹�B����դTѱ�u� ��J	.��� cLA�H7�M��B��嵉�IQ=a�nr��,�H$^D6�.�	��Pf��h�y������z=�:w��S;�w�~,N䱉�^_AQ1}D޷8D�þ�60,S�4��~���R^!E%� _���C�7��o�ܤ�b�Wq�����U^� Y �,�ￖ�9]��
�A�˧�@O ��D�&r��9����p��;���n������X\��8����@��燐N��=��@�zďZ�J�[�A|n�HN\���@��8���I,>O���vJ&Z�X�I��=��7/�(9��'o�gN�׍%�Q�G�_]���uT�~|�'���Ϗ\^^��bv6�勛��w����HiY��J���*��PAK aA	�cJ�����(�� �$���2$�/�`H�緵���L�X~=�	���; ����ē�c�8.+_���9�G�&[ȣ�S�h���m��׋�x)�����.��UN<o`p�LZ96	oD���̜�;��{u����v�.UI�!v9�A�����D�,7x\�Y��2� ���f3[�ǪD�{x����_�����>#����/A\�����.���O �"E/��ˍ���*�W_{�GT���f(�������:cJ<��֪e+$�,�ZD��.�Ӊ�Nz�qq����0����%;c<�O-@�~e�c���=���A�]Ψ9��M�n���{e��p�&7�����>��U����~�j����%z��].=;۬�L�*AԾ�s2S�����~��9�awʉ?G��"??'��ѷ��X�]�-���_A��o3��W�.e)		��W|kC&���m���f��xr>]|Xă��=��2ŬO���+ǰ�L�RT-�e����	��lN�e<q�SSS{���e����
s�����7�L�jtt���.�;d�7U�U���}}$	�G�+��2�K�['r3b9�o�Æ�v=?�AG��]�+_Z�wAإJ@!�>�@�|�y���?S�9���L�s/%]ќH�B�-���"��0�\�t�h�%�'xb�_�j\����~Kl���:Jء�n����b���ڻ�?����~ ���;�d@�O�5�D��Ӊ��b��H��N����?:��Q��(J���0��LU���S� 
��=ٹSd��qJճZe2
xQ O�A]���v�M�)\C��G8$<��Ǻ~V..���Ο�C�LU�nTs3��b��F	�b/�yq0��Zfg���y�m)�EQ�Pޓ�I#��H ��V����\�ƈ�����v\ ���np�����ˮ7O܄���kik�QMOO�R���]�ʲ���w9 M�a����w��������3Rѧ����a�<��@��G���R>v�$1�+���g�^�]�D���S��}��
��(�\��Q�������&i���O8 §N.ܝ�V�zl�]E�Lx?S!-:y�.��P�9���(�G3�=.1ymaȂ2QQ�̄��>���!���rڪ]��W���BΒ?HѶB/*�h�!i��"�Яy��FSW������24���%u�#IC�\������I/vp��T�p��-���}A���soh�'�ӗ���_��59������z#�[�P���1�y�)��^a�=ӯ�v�G�ѐ�:���yP���i�b��{��ə7 ޘ(U ����;��ݢ��$���m���p���OSN��Dm!M8ddc���]�#i��c�[��aW����f*���r܋\{�O���SUK#��&G��9G�	080/�R��0�vpAEy�B�3l������Pu��/���WS�+�ej��]�`Q\�X*֊�	0B侇�s��L��s-����,������ /M~w�>�^��i��ݕ��t9 M�de�]T[XXp P}S��	٠��r���G��O	cd;��&7�г� �7и�(�u�_ʌ�v��ĳ�fnm��n�H��.�<宒��L~��;��������A�'\�W冭n/�7�$ဨ�񃀑 3Y�=�*Afe�>T�+�����bx<�s��ȶ����HICt�r��� �\|�kb3|ťh��m\�����WXI��
�.A�A�K��1��j:�Ԩ^Y<!R�*�C[�S�4ih�6��@��|�܀L��}bUz���!c�W���I[\�V��M�K�j�|�h�oA�>�L�����)靁 �Sc ���#�>����2y�3�;/�;�v&�]��)^ZڅMW���I��<~{2�i��,ysU�1�+� =��v���QG`�ķTu�G6��uf�b�@�M>��Y�2�疵�3��A���J�Gq$��YS�]�j�]��J5h ^��d���\Cp��)Ň�E���.�@	��%|r�l1&�N��Ï�B-�?J�.�m4-ol$â�3R�q��{Ϥv:m�����b�,�mX����\�PA I��K�d��`�%޸�U��6�`������F�쫵��n#Z�#���|tZ�BS�S�T��Z�l�}F���׮�dac�s+��o~��z�5�j�L�A������?�,��rkl0ᾙ�OʢQt�p4���۫&"_pƘ>�atlYE��Fg���Fլ����,|���\h�S���fI��k\W�����/�7��P�N�)��`p�����0ɂ�lB�U\m��������ؘ�+�p�>_��9�)��	�K��)A��(��d��_ul0ZR�K�X����7'I1��Dk�S�zK�?.�V��9;t
}3�<Dk��*��t�J($��X��%'*���m$
�N����.@|w�b^ �omi�����s1T&����y���3�!��I^n�0k\�uX���`:??7m�䒣s�����G�J���E�0T�5�J��nRM�w��8�����������ձ\��i��U���Ao/����JIF5�-B����.��q�zÂ����%ݺ����ِ�t a�ĩL�o��o���� _�½!��2)��������᎒�(�vL)���Gi���r�[�������������������������	���6Ϸ:::�K�l�Th��Ri�Ir����bœ��1�����Qs]�Y�8%���<�߰���qPJ�(%9u^��y��\y��S1�)�'Ա�8��q�}�r��$�L ?= ���T#ן�J�<D9l)	H�i�oArf��t�\�K���
��X'����~gN����f�vT�������͝WZ*��*)O#�3ʻ�7�G��ZDD��Ieǅ�`���6~�<`K������L��N2�hs�I�?������	}�&���1F�u�t�(��B�x��0���J��r��0�,���K�K�.�������|�ikm����ؐ݌/�
��%�6�]��kE�4�Mn5"�Q��;x�(�pVT����"����p��j.�ـ�I\����E��L��F�k��o0WO^>��F�H^��#y��cj�c;:==���Y����\���l�w~�%'?���E�FEú4D�I�w��Z�/.�,9�$�+M��ҁ S<A-�Oq-�1���(
Ó��T�@�	����#/���Dc0��S�����uGlׅx�B�xm`�'��O�-zP����H���^O�A��g�j�,�Ᾱ�y�q��_t6�u?�������/ZX/)�|��]·܌��㝚o0�*x�85[MB��	C��5t}�}�^��E���C��R�����gx��۔�S$�vke��U�pÜiH�/�p��滴	gW\շ�d�t�Jqr�|����C�8�ˢ�{�+��9�Avm��ܼ����R蓉�h��]t���w�G��V������ �#YF�C�}��շ�9?t��m�p�u����)���ȱ�}��?�ތ��Ye1N�����t��r����Ȉ��ac1$�nD�C������n�dp��}@o�ˀ�3bi�l�f�:�O�'�[�Q#l�Y)��3��Z����fU�=��c�v9�M9�c��3G�)��n�� ���GIR]���C���Ӄq&��5,ދi����nh�0f��ix�F�M�lɕ__���>�rI죲�z�Df�%W��Y�퍩�@ <rMK~@>9yh>3&g��̓_�v������G� ��K�,<|;䀒]�{|�k&B ~�
Md0[��_�_O+h0�L̹�� ߅c�+���p���c��Z�}Me�⃛@�O0�3�~��4�C,�׿�䦶���c����]�~!@�3NK�X���J��)�_	y�!)��Ī1��W~���/Ȟ� ����V���j/0w�������*g�]�:��!�'�g�f
D�O��@)~������ҙ\Z�U�Y����Y8&���U7���@+*x�ٵ��
Zp��v=n�������z��\���Qe�^��j�FFF��M�� ���Us6M���ʚ�i�Ӹc|���63��s?t�|}|W�.#�sێ?���)k�..8G���X�G�c�[�{��v|���������F)"B���ji9��*�R�^�i�D��f3��KȮ��MMMʹ�%d`p�`D~@�|(s��+s�tY�!U�SK�,	�JB.M�^�1/\ɲI(V����d��:Æ��ga�pʭ���xm>@"UU9x�
��lTҧ���@ Z����066��v!{sjEW���������/������5սXRr�F)+; ���m���o+�t3��J�b ������H��0|��ȓ�R`b�0j.?{��^RQ1��L9��/�u���!��駵	ؤ�pl{&�[A�ӟd��JM��z����{��f�-�/��6&���5�=l\��>�ᑭ�k׌CLl��ğ�_:�k`@�vA- �������N(XvD6-��?�&v�+����G{Ͻ������,�w��KN���nnnK+�@���zWW�l��v�8��Xh�uh]�*�2�"qܙ�LNI1�727G�k�&u�2���jY��!���)hS���߮,�%��p%��J�:�;��������R�κ�hV�v�1�1�ې{��`��7-�Q�R�a.)���)-m���w��ܔ-��]��>[JTmd"���[&��ʊ��̻��.�bE�k�#��0�#���8�����U�X`9�7U�E������f�I:��~�Yޒ�lb�iT���T�%W��]t=q%��ף]��$e��E�rL��ih����d���}*I��[]]�,b����j__S���7��}��'y�Ғ�䗕Y����O	�G�jz/0h�Kݢ�w�n&�l;M��~���[�8�[�f��ʋ�#�ذ�?�xy%w4�t>��A�*���� a����'|ԲϚ�l�;�-�_�F�s��f�R�P-��-%�7d	�̈́�Bƙ�(i!�;I��="��m��8и6��(�h@s�`EV�"+���)��mg���p%�k��r*}���
�J���;<䆛�i�M� ��~��O"ek�{�4����qQ���
s0�(ÞF0�A---�1�\i��{MY?EC�b��ݾ�?����3痗t�ud�S+��}j���\h0��>�����_6�C�໿�1<u&$$, #�P�����ֶ_�wQ�{t���X~I��qi���, �#��;�I1��}��y*!4n�0Ѯ\����ͯ��&*���PC�goo���頦��S7ڴ,i))�O\��@���Ҳ`�.�$F����띹�����{��dzlC�_��s�&.����Mq�jCb���	�\[�"�9�R���ӵ��&���2W/ߡ5'mr(( ;��K,��y{��g�cm��6;����)L3��~���k{^��E;��J2T�#��Կ`H�$"�^��vGp��ow
V�F��1�j���_���nT)o��3 �'w��C?��].��	p:���+z�������3�#��������"�	�i��v� ݠ���s-�:�sq_�L3T:{C���_m��3TӶ��40����6�� \@d$��{~Gy&���C��{Se��4O%����#�?�`��}��f*f�!:I�Z�}���鸊�摑��<ZT��G@ �6;��2?��i�M��kl\%�X>6d�l���t�8"+ЩjX��/ �V�)�\��q�o�o&{Δ��h��N����_v��<?���׿�i�<�M6�;���;�\NX��_��PٳZ�[��hJ�M�e�¦
7�;�2vh흰#�L�K8tJJ�]M0�{���Od���u���e����dƄquqYI�ȑݿa&@ H�OL[~>�B���o��B�!��8��e����h�J���)�N��K�灶���StT4���:��aj��9!��*�6�{	Aw�32H`D_c���9��:���j\�l:5W����(�N��n��qGGG�����+�B�b{' g��3��a��#�^�B�����@��o>�ЃζF�*�x2�xE����=�#�����x} ơY��,���uV|��	嵔
���6�NA��N�?�gy�������i� ξ0���eA�v�����W�O��/xQV��A���>"�=p:��
	��y�)?�(ι鮭��C����!����3�~�X����֯���רڽD&R3�hMI��>�»�y��v�o�9�V'�ҔeD�|���4�&K���3�l>�nGwG?��ĸHa�� �O�� ��־7B�s"�1�,R�"�G�77��F�B>���4�����fx��� I���&w����`�_k�gj�۽�tFPPw���`��Ǐ��_���|}}��)�����o���>�V��3�Q����.�?U���q�R99�Ţ�M�6�%P�n�+����,--�N��![�N�?�ᶺ�t>��񅆅�` ��ͨ��{��i�{PaЦgsɡȎ����z#�&+e�L�ˤ��F����۱���ܥ���_���8��J͈��+�6�����O�����un���G;���<���0�)��U'ſ�"���n,�xA�h���P$�i����b�SC�]d���V��qP$��9l�;Ƞ�Iæ?��O��p����rr%�������^a�t��BGZ�N��^��L��f:.��e���0��L%lC�J@1�Vj��Nuai�Z^n��܎w�!���Κ�?0Z�u�@�.���.���g!R�3Qǝ�Ke:,��5^:��$��(�Q��F؆O�3����l]G��oyV�[ZH�� nN�`-��\lu/���'�f�I���Z����������N�7}���B��R)��s�t��#��v]b����N,?�����c�:�g0�%0��Gb�u�п�ͭ~��ը�L�S9C|���pv��Q}\�\Pw��]`A�wS48�giJ:M�b'�N_#�׷ۂ�1��L��U���� ���g�u�Lf���Ps�#C���n�BLlƙ��[��P��g�zs&��z�Y�[#�H���B*ŨF��Q�|�c;We�r���DO�Cy��x3H#+������AЎTT\L)�t�5Hԛʢ�0��8��<)�`���Z=:Y\RR0���jR�� ��ړ�U����Z�sK��`�x�!Z��ëI�Sv�uz��rp���J0�X�W���WVQ���� �-̆SPZ�V^^�Ns�1�l` ��O�*A
�M��b�}�ƈ�^�����ӏ�Ŀ&J�䇼
/�E�L%@Ps��4~VBP�pu�����3���Rl��u���]���r��0E?�m�JǑc%4mo�r�}3��^��e�A�[�E�+��W�#̼����J�d~�k��/��������H�X� P=r s0�yUU�ִ)������ɨ	��9wT����]GHII)�&�y=AE�!�ٚ/'�"d�P�[��n���vZ�0�0]�)^e��}�hAA�5tY^����1�wU�����ZX�pq�����|�k;�*ho�����fNV|4�T	��B'��ZS<`�u�Q�x�t�&�+�4ц�x\#��/����^��zкR�d^s3ߪ�����3G���,�Zr"$(d����xe����5���^�݊S3n���Am+&�[sM�19"�}�� �!���e�/�C���Zx�/����М��ta܇1��{������ �CCyH����;lH8-2q��u��
���[m)]b�)���Q����M ���#P2�#Q�wك68��D�ϥ���*	���_C�д���[j �y_WW�5/�x�@dR��b��� �}_y�R�OG8=tt,LL����כ����I���p$���i�a#���P^!���Ғ� ��_�2��`^�А&�-f�ｽ.��+筕�T��-MbM�L���KY[3�2w�H�A�ϕf'ҫ;�� ��M��l�wo ����o}�Z�X�G�tv
z���H��ʀ�O4�h��T�� ҌG%�r*c�ܼ��RRRo��GG�Vj\�z�ׇ`n�6�n�`�k����, h[T�xlqNk��g�����{�4���!wB��y�!�0R~�Fy�}@`(q��G���3A�lNK�����Lhh��g}�đ_�S�11��?WR5�i=??�,WD�:�uO9��;��D��a��:�̹H�O��!��H�b`��H��(�@lu�Ȳ꛷�kk�K���ͻy:�ㆇe�45-�[�9���޼��g��q��r�.����������$����w�W�<�_�*��
ev�0����b�'��� e<�[��w�ᠷu���`@����@����\baV�lmYܠ�R3�%��#ha��ֺ/�������	^�G!��	Y�l����D�;~�_�i��\�#���� ��qeM�q�Ր-�K��ph�>�T���v��p"D�����e���}1�*zm59�@X [��AS(Xm���J���*�.��tl��]�5�n;͗x��y	Ŀ<`l��#�e) G;�2!=8�D�0�8ർ����q�ߎ�p^�R:�T�����d�x���h�kE:pa���L��q��� ~z���D��'*�?��ħ'CJ;s�O����َ�ڈ�J�m5�I\~�k����Y�&�<�q����VT�,
�h���[�Ǝ�!��ss��\o[��u.����2�һ�P2��ޜ%�7!�+ �����GW�KjqM��6A��^o�|)Y`m�i
�a�L����V�M�0 i������X��{�0�K M�LsqEN��l?�9y�����n&wn[�@��
�wKa �������V��O#��\���4�leV;������<�D�����y�F�[6QYS3���q�>
V>l�C�N�����Q��Dr��i��7yqԂoë�;�����z,,,��a����l�g�^%� ����GG��z7�J�����r�/H5��QM0�Zɀ駪�:�!�;�708�D��4^�,�K�J�i>���J����+ʹ�3��3��KM.�������hZ�0��/Y���zvzG���Hچ����ԟHql'>���ڒ���^^^�a�ܳJ�����ӗR*������zuQ'�W|�3�wU&:_�%^����|�vT��.�;m ��a��_��er)g�nnnZ�ۇ-�rv����e��l"���m��^ER��(�$�(���jG���hY�Tn8��B7�w��]z����Λ��t,@����Ay��·i3k�ɟg�Э�f�~ �e�d��,Qy���.�e���n�Ly0@��]��:�Ȫ�:%.Z`��t��&щ3M/(�b���1��;)����E�d�D��e��F�V��{`~�̈��G��f��s���_�*#�q�n�m/����lbܦ�iAT��y~yG\��]R���\���5� �;�ٿ�o��� :�fhiҰWf��K�vvf�ZP�kb8��vH>�]��0��4l��-=�HNM��T�<K��p�3��i7�S��1~�w�[��`�cx�0��"��>C���-��U����QM|���4�WB��~I"gM�;��n\�S�~����
�8�����m��\��C� !H������-x���{��5����������֚E��g���ޟTUW�����-;44PSS3q0�t��:jv�Ò����r�1؆���I�oi3��Ʋ !�Z�2"8��>hll,hg�����p���G�����Z�AQ����Ϸ�T<8��}�P�1=��&(x��r�{�u�MC�>Q���)����XYm}�e��״��`� ����l=�H��m�7{��_bp��C�A��x� �tS�׍b?r��5V���-�Z_(�Z#�}�5��9�$M��h>�+�L�)yN]���l~$�YmT��T��+հ1?@p��
o�g��M�
O���|������s������QdT���~����ݐ�g�=BL�.�~}�C�Ռͫ��0Ǡ̌�͕����rK3�66J� �
��cM\�Q�,G�oH>Ȑ#���#e�D��̬ۨ���@�Ȅ�q=�5P�!�)�p���8�;�6�k�!�oM���r��$54p���S|�ڛ�����f�SH1�:D{ �[�t��Y��u���Q�e����c�����vij+�Cc�wT>�bi�VZ*5}��;�C�RI�!S���_,��𚆧��4�@��UȠ�����*�l E:ͯ�aŃ�u��ʴ`�蠸���m���ƒj�����qg͉���0"�g%�S��?E�ި�2i!��Tٮ
/9��~��S��ښ��8�Dc�_4�w�E�4�A��+ǃ�g�ப�an�;�L�$��d��r����+H/֢m�.'�$��	dn��ݽ������v�����XT �P�A�r��}�֯ϴ
bk��*���*GT� E��ߐ�~5�i?O��������r�0c�tȞ/@<�RR���0O�9}�����|��#J�ғ�+�TP+�z���)M>���T�}���#i����_s$��Z�i �d�uT7�-E &�m?�"�V����(�?<�~�|��mp�%<�^��^x'� c�C�|KY����>&
B��Lq�Kʤ����#�/�����Y�9�4Quuu�22T�G
�߾��5Z\L��@;�m���-��I�+""�$*��B z��Lq`���냺�7����&�2O?�p����L����o%I�:I��Â�"�Gl{�+3��i��CzPQQ�u�E����*Z����&���Ĝ�8����\/G�'�0{�����y͔�D��a�	���T��}������_����a��<����H37 Juk��.gזe�ۻس�+ͪ4!4v�PǸ3������.T5ӟ\会,	���v�V	�rܯlǦ�������h�G�ϳE*5_.���Z����� ��u��hB��3���?� ��k5����*��?d����L�Ĉ��Wu�S̻�>(�/=T�pM���T ��\^��j��{��Nvmj~K��~���~b[]��ݰ�#�����fN\���I�6a%���UQ��k�ֲ �j�o~�{߄����1�ɫ$J	�%vy�J���i2�tu�QT�������o�]7�uv���s�r���gl�������]�����xb�珨���:�ٝO3<~z$^a�Rmil�n�1�Ǚ�u�c�e"-m�G���	�⧻�l��U�5s}�fk�9�� ��~�8�����Si��F577�D�Y�	�߽�0�덭*��t��_�*����S��C5���bRܥ0!���Fi<:���9�����+�1��2��͢dj|��)ͤf���l�f Gd��r�>����L�F��'o~g�=[�c�I���!�zx���п��^[_'����XxHϵ����2���ľo���ZҺ����m߿O��Rݾ�c̺\U�вg�����|jHf� ���ed*�ǺjQ]���'�q*��`��RQ�#d����p���#��# ��ZZ����muF9��P4���YX�MLh�N��u�YYY��_o4�لS&E�^)p0�l����N�ò��8��S�kd��d��}{���쵁���*�u���F���Ʃ�;2�#`B?7w
N���QS	))8@#:R���|i�Q��o�|�)�O�~u�_Ad�x'��`�r�Ntr"lY��L�(7@�b�"Rh})�C���FDn,����ov��w�|p�ܲ�.:��?�"9��a!5��=�������<����U�o���m�M&�zeee*0���,�,��]ʊ�xQ�#���Br�x�_罦f�,uB������R���G���='CCCʽ��l���H;��!�4 ?W{佉;T����>�l�m����Bmm�ݖ
��Q�Jݽn����ۊ{ɮ�o=�� �O�Q��u��6$�v���o���xI~,EҺ�Cv�\^�njj
Z��<�Wڽy�����5?�U�� ��yF�膑V�;��\�Y����7^����~qt����kY�Oՙ���+H���"Z�`H�2�MHL� ��楖X��*��5a���Y�0L@�c��.�YP�x����\�D�֯��|F��|�(�U9�o�f]R�pg-�M�~ �1��!PYl�������}°kj���� ��ų+I�`L�8��C�5��f���c��t����g@(��ңM/���uI�������R��H ����M2Nv��}�ڌƧ��ϣ���ʫ�@����"}������2���ީ
i�´�a|�=�Z� 9���oafX9d��LI,����f;�K�����ǛM���*{q�9 =���xnoh�s����QS���D¢�"zF��R���H�U�iEm\���O��G?f됿;���$�xY��b~O:i�AG���|ú��{���4�x�Ȼ��q��U�0.A��Nm���}}}��=sɟsé� ena� HU�������}�i�يͱ�l��>�9-н��3�B��w��+	�eb(�{XuA\�v�92��3�0�~Jɢof�t���Y�v<����	�Z��sm1�qT����eͥ��l�(.���ێ�����n��*���T;�b�''gѹ��+�f�gƷ��.��}�frb�GYU5�ʌwO�]����z1*<..�+����o޼�������l%Ad ��Ʃ�U��c�F?��@��}�=���W��|�5=a#�����91�����V�J^r[W�����Mdi=A����'" +����f``���� ��j���x.�V���*���>G���A���{l�X��nǔ�qV�c�t�3|i�S�w<�S��-C�ܲm$G�������5׮�!9�6=�$��:��.}Quu���2LTxv!�h 3�&�L��p21IjiB�i�0K�ަ����/�jO8���R�{�� }����-�e�BS����°�$q3v�BEJ����C݌)α�;Y@:�tGRM�`��p����y�s�5(&�%(urZ�qd�/5�" ���h+�Ã8ν�=��B}�L��8��<	�m���B�wz��f��pr�в��@��[��͛���n 9]\��b���C7d?�83/���E���׸�[.�l���������5)�otD�a%���G�)֪�5�PLY������䉺�k���A ^^]���S�}*����g`��ma��	�2*&@oCu���9������X�\\���u���� �Е�K��������'q۟M��[�� �J鈙{`�؞�|�eP�~�!`�{j&$�B>������ 7��*V�|����^�e�1Z	��d@)�B*�
7�z�ܪΙ9
�Y, ����cb�++1"�{�[U��*���P%��Qi�[���7`4��9���<���F���5���똣}K#C�M��v Ͳ&7j���fc༿�l�?]�="��9Ʃw��pjՔ��Rn�,���:+�=o��OmװҹȶM'�Rb��'�)�IZ#ү�6��;�b�蝦;�؁'Qi�Ln���^�n�x�J � )���X�85А�����~{�:�ħvP�*g��>�p�&q�jz�t��Q�r�54���+�3��tY�@)1;mv��ۑ�9���%%�||��})(*~w{%�*ή�}�\l���͏�V||H�����oSY(H��|��M�=��]���z�v���RfP���ņT*�"�qܷ�oqyݶ4:mU��z#������v��~����H(���[Ι����,�[/����;�a��u�*�w�ށ2GC��M�Ӂ�ZY�SPVfm���Yy|�`$;}�����#퐸�p� ��6��/���K��dr�f=���J��8�d0f�v�Fd�:��ߤ�yw�<��Z*���-��<����F���_)�����q�Cߨ��i�g�c �J�p���?I�,E��xc��Ν�"wHRb)�%�DSL�G(��9�h;��B�>����1��$�xxy?~�u�:���T`���ݥo]�i6!�~[�ef���)2$j6�W�����'?�"�����\�6 �q��:�|�Ց?���	�S���J21��ƒm��JpXR-�;|:|�DH��Q	�+��h2�omo��h~��؊��OY�����wL�%q+�E�լ�WM-Ä�o��ڛڡ�G���.��Mϓ��_6Cٞ%nCY}�ȟ'B'��k�s���I���Cy��٘��ʇ�@k�+\�ͳΝ������
LD�R� ��
IQ�M:�{{b���溿z��^HCD�`�]h��ma9�e�E�Zd"��:����Q;$	�?�LW%�PN����'D/�u�ۦ�nf�AY�-u���\#+���b%)!��m�B�k&�!&�o\�b��g!���屍uSȶ�PJ�ׄ�āS{�jj8�P/eT�����<@w	�Zȵ��T�: ��.�z�s)�w/
��h�4HO@m]��%S.�2�s�UUU4�"bF�>{e=at�y�\��Q��~���q4vpy�>��J3!N�������nJ�&���⾾"�.-�c�Q���,e|$�=Wc/�tH��A� �+z��T�W���F�KMG��8s���Jt����2R�<=	��L�#Þ��؆� ��2�f�j�c~��`�{���ze}�j�Bz�v:n��k�}���s�wvv���p����9�WA%Ij.9�y�jl9K�62;*�^z���r�n��pἽ������IQ�X�����x�`#�[?��~�?�2K�s���d����`���ĶY�È���:۞���i/�6|ꋓ����Tj|������×] i �/)@ġ���z�P ƚY]NB���6�H_߽E^Mg����|oHw~� Bh�?1��p!)r���������&<)(#�g�gO�:��M-��^Cv%��m�U�_K�b_�����`A
%�C�X
yx��d1���uﻎ�F�ZY�ߏ��	ԧP�� j�M� �����v��W��A�<CD�ߐ�nl�w�tnsG6[�d�ʹWJ�i�Dx큁�����+�;l��^k4����������
c��d̫uҹ���#�ӑ��_Eo_��4�4H�NMM��ZLXk��/���ļǅ����eϥ��������ݣ#���i���?���~Ki���c���Q�H�㋀O��廪�~\�Ý���^�� <͸ �X�
$xcz*8�%@y�:a}�433#�y, ��p�"���nx�7��Bw��q��so�{�<?=�$�(f�= T��|�ř��������9�&Y�);?wz��?�#����u	�Ə��y�KHo��H��v���V��v�(֯y+8��lhk��~C�f��R��^>��FrQ6u�GM9����8۽������NTT5ZC���A�n�e�8��#Ԑ������!��x�{4
)}�	���R�!s[�Ĭ��0Y,B�rn���;���:��d�v��!cq=��Ǘ(������	j 	Cɕ�u�xvQH�M ��/]���DJ�+���C��e,���� FӘưj>W���n��6l�����G"���Y�T�lr>��4] 8��$�Т�����n�V!2X}s���8<�F3�&�lu�t�u2��@���}Ȇlk7����Ϭ�HCm����0Ʉ��ev2W�*9*ܳPv�Ug*.1�Ŕ.���5y'Hc�FP�gG&�r�=2ĥvg�R6�{�M�V��1Q}��ʢ��B ���͋�ӓ�l֏�]=-��D�"縋�T1��Pl$���C��[�*ZN��6[b��JrsN��>�M��ٵ���{ N�FxTl,k[;y�t�� U���Ⳣ�-ch�Wy'��LP�+_\��ZӤ�c�.%�ܜee��)Ťs�[��9@�f-�^kK$e�6�U?��G��&%`�������D��!��Ʃ�x&ͪq�D�W8��0c�v��f�r�r�Ѥ��~��v��T	;��&t�������Z�Z�e9�f+�49�u��H4���eZ�6j�5�.������Gpt��
oἏ��zB�[�W#roܞ�&��|NNN>�t�:�����J+�Å���۹�e�멹������)7ph��0�-gʴx�g�F���Z��"Q'B�8S�&�|mNC�v��#lrrR��6B�������N���`Շ+����6�L[��i�D�S:ߩR�_�#�4�j2�^���y���{B�@��'��/�kMz q�1t��	�u��竌f ���/���)5_nÊ#ɡ�_6��I����#"����ɸ���J�lƸ�浇��nI�X������{�%Y����K�d�����g�x�&f����.�v(~�e��4%���,�@vT����x��}]@^\����{r"�*N��aww.c":��|6po��}εu��� ([o�u"'��X}r8K�1��<u����~�:�]�|yd��M��g426��1��L�(�\��é���{����Q֝�Q�S��o����s�ٞYc1���@;5 _)S��WGZ �����W7�ϻNo��9��d�=��l]X�R 9�A�@�+�t*�R6#�s�sh:�%
�v#_��@=�ʓ�<^2HR�=HQbAV!�<�>2�S�s�o+��\���냀tC���1�fl.T�풄�hv`,�Ւ5� ]���?��7K�V�~��κxܷ����8�I�K���	LD�]�h]Q��=�-��=��˽���c�s/��KB��C���g���?4
J��c��"�o9vƂX�%�>�ޜ�'�=>������DKC~��A�a�0H4A����l���l���#=Qc1TGn��%���~cV�U^0�i����o��x&ͼ�{� ғ����t�Jғe;9U2����'��,x���	�`J8�xqmAR���NPKr��ײ���h}�Pbp��\�������*dGe9׫�'.����		}7�_0jXĊ��J��g[_7 ҹ��n5^.�͇u�9|A��X}�h�3�+f|]d�D4�ߙ���'��z��om;1���oH���X+��"����;U A+�u�%�����. �$w��-3�5�'(��=H3���^�R*�����
���f�:k�G���/j��d}ʾ�SA���y�����i ݠ�������#� \^]1{f'��Fw@�*N�w�~�KkZ�]w��p���@���C��C�a&>(_�����>7:�d���ȵ�@��^cK����K���,���;	��Y�W��$x�����9�����3o�F�Ԟ0U3�x
���9��&��k���F�2r��}(x��vJ�I@҂|_7�$�Y8��P�N��;�n�C@�n��L�\��m:�@݃�����&��ӓBH�Jr�7�$��l\\A���n�947�Dȧ��܂ܪ�����
FQ]�fEׯ�C�������IE߅i\�o<��*Q� 8��D��R�Ѷ1X�.�>��s��PbtK�[<�FU����@���.ϋO:��F�R�l�� �|�c��9H
�6��r3I�Q��*x� {����.v�jj��"c �����3�q�B����2h���s�n�#��P�!ЃU�FA��[=����[J\2�|+$�J��9{2*L:���B��O���B��KjC;�zρW���	ߓHזp`�>�!�Ѯ2���X泻W����u����R/�����7IO�ȯ��'ޖw��d��}{���G��8�6@��!TĢ��H$�~��S���sBb���l%�BJ�8rWjK��:�Q��pZE�� ��'��Ԏ���m���o��Q�r���ң(Hq@ۧ���%���C���$À���X]�0F0��D9�y�:p*��1��@�F���hq\`�!P1O��*�椠���Sj?��קp��xR]�/��i
�Bk�1�%����rTPV�����ϟ?)K/�Mn���:�>i��4t�!�wQj��O@���1~k��;��Q���y/�����&;3���gLx�!�P=!@�Q�QY.���ZX>�6��:o�N��AƖguH��M�ߠ��p��CyB�@~����Y�_�&�zr��۸'�;�}q舦��zt
�:�@�&1@�?����w���^�H?�!X�Q�p�'�-�+������p&\ �@|�ME�\Ջ0r��Eh���s5D�l����:VV�����Vip/��t��v7�r��y���	Z��74X�/'}��YW%�@r�
��0+��w_l�Z��O]��7a,��bH�$'p㓬��|�j"ݣ�$�7�̋�:�s���xxx &ym.��$$�rP�Gvm;t�9s�'��U�+�{5yNE��� �Tj��c���Pל�*\�1���� ��]>�<�k�t�yxV��k���_��`�����'�ߗvoۏ�|�@��-B��A(@��y����ls��l)�z׼F�[���&�I'����%S����?�A����fB�cBp�4�zF.0�Ho�]��/;:2GM�� ���2�&&���5�9�ʴ�V]�
a�����O}�R<]x���J/��ȴ���G{4J.���<!��;�{gvr�Y�ͱ��W����A'xs_�����Q��/���p#Ĩb%l��m:V��R���u�e���!<�?�&7��~T!S�Svٟ�z��R|P'����A�>�}��ˏؤ'#J��ʔ�K���]WnE8-����.h阾���2W�E-mF�V��Dè��d�rm[��x3#6�#H�X�P����0U{
S���%�f���)�z\J|�@�F��B�2����1z|\h��9N�R*k.- �!�#��a$2����s Y!�G{��2���t�rs�Wεx!x�uO����l�F�<Y�+Qb�m������N(D��춺+�a�y̲�����9j�f/)M�L���-%#)
��A�,)#��O�G�=e|�]ZQV#xB>�ǟP�Z�1���[��������:s#(3�^:� �����h�Ԏ�;�۲U��-�nD���UZ;_s��ŧ0帻�c���=_w�o���<�����sʘ����Oϙ9�Y�؉����K1ضs�>:%��X������d���5��٧�8]������@��8/���K�r<�����WN��y�����>���q����/u�M�JX����#bG���0"�ow�0#	X���c6����Z���,5���n��O�iF�y�@,��iӉ�V�!���w��$c�k��L�3K��c��t�ي�F66����k���|���}G �T��Q��"�7D"+�"�,6 R����U}?��q�����[��oé�l/�hWY@a�p�݇@�<\w�Y�"ԗ��*6���3���7
�;e�ڮb�m��0�7a�o;5NZ/�^�^���h�/À��(��<�8�~���4\��B�Bz\W�н�n9i_�(T�k:��hk״O:E����t=�~�	����	FZ����iNEh'�V;m�_��j�w�
�P^^�z���|���@�:��v�U��v�]ߥ�+Ъ%��b��	{�����9��<����nM<�}~�=�D�%%����e�0�%V�����Nkr[�G|�Y/۞w�B���7�����&�����(�T��8|OR�9��~UmM,C�U^����ol��mn��
V�n�d���*<�
�%J�h�)}��'f��{�� l���D�a��;�#��%7�~�ngj���vv����`������ͼ6%���*���s,$�v���-���ڸ��`|�=Я���o��]�l+�������>7%~�f�a��R�q)nl�����q-}�ef�����m^Œ_�4HP��	���^v]}b���/�[�-JB�"�{r��r]��c���Gf`<Ht뺅B۬\�C7s�B�AF��U����*Ha�cq���ܚ��'���ˍY������/	��U�vO`����x]s�[ܕ�D��r/��KK�9323�ݵ��H���^ƚtЁ� �K�[�9�G-�az�F(��2�/R8au,��g��>��u��n0��5^��	��h��ֳ�GM:��.G��g�й��,�E�~�����U��lSn	UKE$��I\P�g�e���+�s}x1��U��iで+�L�5g4T�n�G}R�ͤ��Ud*�r�~�߁2�����U.��XZ	�z>���Ru� yG�Ą/��#����ؽ�^tad����gi��[��ۍ�(vߕTOl
ؑb8�����ǣ��O�-�ڕ�_9�OGC\�_tB^�o^��_![g�>cvЊvq�7z�gM��J\��Z�AN�=������-.YK�ZV1�G���;w4<��?�9��i��#�bo��	�°g>i��_�-��w2y����t4�@#�'m����H��s�>�E,Y�S�L��K�J��*�c ��D>3T_��***�
��W8�c`2)޳"�@���n��-�Md�������Y1&��̌������g�͖B��;���n��:M�o&�>�sp(�~��@
�����_�z.y�{ Y�X�	�䠲�њ����FY���FՒ;A��#2�J���Mda����5�w7��5�$000�GGR���:��nή�F�?��Qf@�Q;���OU�����{bƱ'�Y��]�|�V���Ό���,��j4	C��?2��*%"$�;s*�a�)�ؗ�G�>��	��e�C\��R�s�=�RI(P�]N�z˽m��_5����D����:�>/�uf?��{BQ�����E-a<�6��>��?�?��u|�9Z����=a_}���}% ��^��>#�f@���%�1�3�rv���QXQ�,$��fe@^�W1{�>5Hcٹ�BT���P!;p�3 �i\�V��"=��P:�3IT#D\\\_**Ї��)Y��D|k_l~[���


Ԑ�����"H]b���e>gp�"P�d3��mF]S�z���Y�U��gE.kNA��+�v����ZV&Α.I�v�(e���BDDMR<e�� �p```�pi��
��o-�o��Ym-/�V" ��:�����X�'�O�J�F����Eb&+����/A&�����**��31)L��CH��w2x�ɩ����v�#��؎ε!�җ%v$�HI,k]h��Ob��� �s��E��S��=R���ԯ7�R����������\�x7�cE_�^E�߾��������y�F��o���
��I0	��6j *�Ϭ��ef#���ׇM[����p�SL�C�2�u�m��>z���#r��c���T�y��29�nb��+H���A��in柞���G�#�*L�`p�LJ�7?���e���UӉ�1Ϟ��R����]c�BY���,	�f㼺`�dm��Ey\ұ����]�gXpQ��E0fX�!�������Mk�8�ƒ|��L8Q�� v�xд�_�?��fQ�3�m���<���LJ�;�|�1��o �~��5���8/v�z���x\������S��O���L翿��������
b*:;A�xd��Ĵ��nU&����!��w����_���4k�M{&��#}��Cs��x'�p��m�Lyfc�=Yȥ�r��.����[��?Gը����6(��n���9H�$g/Z#YZO���Bߙī~.}�� ��h3i^���i b$�7�kW�.��3~~h�n��R�2��z���1�"wH ���{�¾Y��܀�c�CyfbF��&����-��?~��h�n�AؘB:�58�Ywmu56>�7����8���Ň���hw���e�f�)�]�HX@�x��х�T-�V[̨q{c_=5~y����(�?��,�
�I�þ����ܼ�JG�
\��P�S�(z{&�����,;�h��{;−D(U��=���X��(<�ȳ&}f������ܬ�5#��t/�\ssq)<��)N�����tQ�M�zn����w��Ķ�Y޳��6�T��|��4<'ze!�:2�1��`���4{O�X�= ��}��Tk�c�+��?���[��&DO�W�YD�̽�퍸 �/���Ig����`��:�pu�]�����W�U���Q��Ǯ��4��,d� �	砥�9G��4�x�b�H(h��&���$�^(U���F����y�$I�cPkO��S���s���m8�)�C�^*+1 %L��a�!K��EA2�3E�����p��(��2��y"��	Bp+���-�e�EK^Ș3D��cIR�y ��)��1Kԛ�dŷ׼��*��,\��Y��d�49����E	�.��J��0�����\�`  �7]h8�G�+��W;���	�0Z,�4H]�6[��f-�*�2,��ի�/I���ǆI����$D�έ�c�g�,w�^���Akm%�GrE��׊�U6����ճ�v�t������-++�������x���;������{zz8���*;m�1�<P
�a�]@��l��d����%�|Ez��+p����Zy�r}i�H_C��xK�D�(dX?Wt2(�Ea�P�� �=Cɔ6~wM\+��q@��`n��������w�)�A:߁ȇ���t?#`�}����&���]���<�ô�����Z)W7 ��mF�[yO?D�mEE�QD6��)hi�C)��f,]���;�B�%Bw�y?΃
S��Zl�sێ�@�/K����b�P��I�@U�7f�^�>ex;n�Ȕ�!cS��	4�7�B䇺;pm��Fr��d�ٻ<��3؛_!1Ts�ll��̩B�yZ���5��u/O��ڢ6�*��1��GIRbNyM8/��p����\tLAL����5�~�3�H��ԃY�����z���q�t��)�����+��4�������]���䤖F�o¤K\7�0��43錪��K� ?�B �μ��_�1�?h!�^˶�6��
��.&�����F��Y�ʖ/}o� 	��;��������0��!�()�L׻�߁@t��r��)f��&��ֆMq
�ǻ������so�̂�an(#�������	9)��n��Su�����^k�N��$��'��z�j�S�4u�g\���H��	,�0��HMB���GH9d�j�g�,���ת�3/�1�_�mk�wʼ`�C�TGLC;b����� ��{W��ug��C>��6s���x&۷�Z���ON������"/�1��κn9��%;��5��z|�>%d��XHaI)���6��Yj��������15���Q-@\��J�5X1:x�������L�FAii)����f��~��U�(�9�{��8"%N$;��ѢM:ǽ��9%$�
�3P���UR����_!ߝ"h,�s�4<�d����t����~�����%��%�|��_Q�:��D.���	��:.9v_�_Js��
TF�~�ؠv��L�P�"_D�pjV�0��|H,��Cڜ͎��z�������q���� ?�!�������k��KW8p�ox-W�֦7�{;�8d"G΄�2f��|�k_�Q�毬�o�)�$$\�fnE�ԙ��k�YW���)Z1�k�p�����ي9	�|F\��N�u��*K����ܶ��~�؇��7���h`�	W��ӑ����P�yPq�UFA�->�+C<��u'��ۈG��*V���S2&%��ɚ�NZʆ̉�s�*�����Y�U�L3�����L��_�K���l�0�=��/c�}��˘x���@��ڎ�K��{n/���ᯪ���B6H�'A,�����BA��ߔ�o��r���p���p���śY�,5vΨ��㤘8;;9	�{ �G_Yq?0SH~�t�����L���i�l-�Z��[q@��C�Y9:t�~ӽ�4��М�ן|����ʙ�����/0�u¿����I�J����5$N��p��H A,���A��ɓ6�E�����L�hЦ6��H.��h�ėH�T�arq1ryYhwL�,�"n�R�S�M&с��b8Li��QD��Ks��9�q6��SN�uB˂@��'��5�x�F���6�J,�fc��O1���K$Ss"~0mN��,��5�a4�i�&}��ᦦr.�/Ӿa��i@�g,���yBB#�4[Q(�:�CI>��:�S �G�ӡ$]����F�4�P
�5�蛿�ǉ?|��Jq^���W=�Y�8��"LJ��x���l_�5�2ב�3��z�	!+۱rX�fx����"Q�趸9��[�Z�*�P��ͨx��Ge�PX ���,F�?����3�%R��@º��Y�<#�ka�̴��Vx�V7���;���'��������zV.pA�T��[a�&�5y%�P�la?�pF-V-�����(��	Ϙ�d��e� #Bo=<�:��Gj�����W5tXSH�]m���Ts5�J���}�ރNA���#$b0!���?����g�:ʓ�<=���"7#z�`{K3:ԡ�#�=FS��� 2[5�N�4�.w̅S�q� 0��O��'o�k���:��T�/�9@������5b�n�&@�:��9r��^�:����PPۇ+t��
�y�_�@�:-���m�ZA,�;�5=��+�W)LjB��5&3�X^���w�j�:�l��
�Y-ܝ�����4I��9��-x*+I��B�q���DA��O�?%e�^��v'�a$@v/]�;,�ʯ�J�o�(0�ʃ��5�	��T�����@	ǌcw#��hR���H"W�X,�a����[��Is-�ƊȜ2���Qi�Nv�Ci�W8`�L.V�J�a��	Jvɏ��C޶����f�M�qȫ�,tf��=f��F*�E*Ѩ��������'fgC���[�$}}Eb�.^!�.`E���b�3g�����ˤe$���e��4���S���#�_��"�	[D�NGZ�.�d�Q�H�Y�%�)NNN^bW����뙦���@��H׊s ��.��e��]��!]�j�������OF�Rz��i��$���ϭx����J?�VD���Q�=���W��%� �!��!��1��-��())�t��]A&��IW��3�K�:(<�R���Q��_�_�Uv�~� ��d���Qv{��)N,�{��3Ƶ�u�Z�a���'�k�Zr�z�x+�k����?�o{Q�����Pt03BܘR^���y��cJ�i���H��s��� ?�=�oo,	�aM�oZ��K�v@X��(���e�ۊ;����tk렐Z�9x��C&oVH��#�2�Uيc{Ӌd�*�	��o��|ᠣ�z1�Z 3���>��#Fra*^WK�?+���w���� �)�S4p�vZ�۔q�᚞GԒ��Gܿ�����_�P����l�x-���=Q��	���e��Q��B� (��B�K4Ѫ���'�3��-ݳ����r��(i|��,�|f¨����������B!}���&��!��ϴ�.���	h�3�W���d�d�d��d��@Sww%���CI6�`?Ml�	�K��2�ߛ0���Ɋ�Y�X��.T��)/���eP��#<��1��2��!�W �Z�t��÷T�z��%g��bZkE�o$>7��������)_�Ǒ�+�O;�1^�tZ���[�
��N1�9U~
�B�0>�<�7Wd �'n4 l������@�4Ux�l�p>���x�H�������P�%���%|�,�5 ��Wc��+*W��>�����bF�>����}�rcK�׭w9Z0{�����H&y�7�-�V�p��pc��m�x8�jy\ޝ��w�d8��L.�s,Ч�~�@h^��4lϕ�a'LP�ճ�}sF��q�5��"�,��c6YR�z��fnja�r%=(3l��B�n�9JVe�q�)�J���m��C�ۦD���쌏��'Y����^ /���u����f]Q��-�+��1J� A��x���?财���1��d��rI���_� �ʹ\��\c��&��8䌬w�G���~���WQ�r������ ��Y-�2 >·��U�*%?���X���P�a��(�/N���&Z��Ac���Y��PEU�R���Oo��T�µ{w*$+�J~� nv�F��Ψ�+D�`�A�	�G�n�)�UQ�ht~˅9�䀋
�t��I���1K՚`�!�`'� Q$���Ϟ�#����<s�[`c�'�Op�&i�	bø��(��(~�VS�X�O��b"�0�%M�K^��ʴ��S��U�>a^_g[В�/��6��D�- ��x�l93�����PA�9l�+)>��z���`����g����[�k
�~օ��S�Cb_�����7"YPF���kcb�h��0[<P�嬉�n'��8����;�/d�c����b�z�NP��ޅ-)�r	��I0��xi����xX��r�s��>m�����ε�$�DD��"�E-J�����;�Q��D�]�6J�ha�т轎6�#������>����{���k���Ȅ{�g5�SÚK|����y�'�no/�遳&J@��*_�:���1�9�v!$_@�����!�J�d@LQ֋�w���� U�i(��r�lx�M��U��p����)�%d��V>���K� �O�;>8�TC��b��\��$��9�������7xy�c��"Q��d5��s��~�A��-N��LN�d �IR���@�NS�'��������ׅ��l���Y_� �?lB��yw�^�2'*5�(�Ց��-����ng~�`��`�p �T�� D�-�,a��"�Rs̉�IV>h��6����*�����!w�[���bx�a�����}r�{z8I�$����
 Ʒ�Va����o�����ϯ�k�䳉ט.f5��9���, !���A ��!�	Oʇ��ĸ;�x�C�h�z	m�]��5܅�G$�� �=ȁ`K�Gu$^6���S�R�Y�E�Y����Kc�����I�t5���L7"�s/�W4r�?P��3�`�qO�f �;�C�?����e�P qH�>ݤ:%���ѷJ>q-}.}�M�j&��r��[�+�-�y1��Q���O/r����L,�|?���
U�;R����q�Μ={0(i��t`t���ߐS&���&���ۍs�oO~�"�� 
A"̀��w������\^G<K�y!�\6� ���&���>8I�~L 兵"�XU�h3A��<��@U����ZV���H0\6��Fdʛ�Sz���񄫣ף�S��9'2�W�^Ú�r�ԥ��u5K_��Z&,�-��������M?�}���?m�S���Y�<%�9����vRki�g�Yw��|Ի��%'!Clxn��~�m0�A
Plp���%�˰}��D�
��oV�Q��H��ER��Ҵu��
��K����{�
�r���%$�]ox� ��\$C�P���1�,�,�R�q��@#h����O�237D�"k?> n�9�x�PXwT��¥��%�����I����~�[�3�q��6%1p~4�[��":1H�K�cL�|,5D&��T8��^G�*�ǟ߈�l���]~.�b��p d��/��w��E���2�|_e�Ȝ�V\�d�`�����g��'0	��Ck
se�j���7���,ֿ�o'*F��W�P�WHѱ̑�޸殭f��N�.�+���H�>��h�s%F�u�	��_�d��+H��?A��^ה! rZ��,�2�(�~��ǿ�3cus��o�T�Ix{��$��r���^+����p��#����呡�1J:��;�\\�H[�{��ب�z��
�ai���%<K|x����7D�㼚���Yo���#�)��U��:�>�ר�򏁐�zd5DV�#�)s��}3���+b�~Ne�35��)�������v��zg����Y��1]�k�{�)���mB5f~|���&��T���#IL�X�mH��l��OV�8bCD��3;����Gt���<�T}���{���yg{�Ckts�~��P�%o��ǎPV����	�%xG�s��NAI�i�e_R��!��4�)Y,v~<k!,��1��ah�ښ��a��ge��������)� ��d�~T �H[����WĹ�SƯ
 b,k���BDpӕh��.鋵�Zkx�C�ޚ`r!L��m����q��ǶFr��^"D[�⌸2x�%WnH~l������Y��{�\��o�J����G�ZJ��\�gɅ<~������UU�h8+.T����}�H(�� "�$�L�n������r�9��+Sׅ�`��Ef)��׭-������>%do��@�x�Fm�s�������/��vnY}�	G�R��pi�r䘂�s��{��g�����?�7�j@�<l�ueN��\w
�������uV���m��a��k�����D�K���&�i�s:�mp�m�A$�T#h����Џ�7���À/��p�&V(U�2� =F|o< uH!�IQ�����k�W�xs����A����=dD>^�,���`�P)J,�}�I�^Gۈ%��	(~Sɞ��0ᴑQCԝƀ8�p�/�tNǖ�����[Kx�:��9�Β�+���u^Ѫ��El�Lq�A��w��`��<�
�,U�8%T�c�8����ӘG�+����%�jM�L�;���t�6���3�---M�U;�u��EyMO9@��v��i�L���������,U臢c�	yI�1�T�����¼��l� R%|�4�4��һ�	R�,|��ܼ�H48��a�����DȬ��vi&���z!�_*R��~�:��H�5�I���0�aJ�	�rΩ�n����h�����y���u�\�Z�D%0�6د�US*0H:�!���4�fn�Cv�����'<�=�L�r̀6V1��uYh�����X�� ґl�Rm��B)�l���q��<���įN̨�V�����|Gl�黀zp=w�u��n��+[�^UO�uIV�U�qR��o+J��O�P��e��y��c�y�l��τ[�Ʋ a��Cϭ�=��e��z.�����ZN��GN�u�o��Nd�ʋ�Su��U\�����U���� ��^ ��ஆff�<�� ��K�UB�/bw5Oϫ�u�$KA�g	�w�TR��`6a�+}���V9r_���
��S$x�;�����ؼ8���8Ċf���$�)7DH�m������.Y6�񽧱LŖ�{�����Q�zW�Uz���0��I���ҹ����i��n�'�DT��c>GIj֓�W��'@J�k�iĉLjp�(���yo���C~�/��H)qh�bp˲���q����L�	Li��U�n�_a��F@��M$���9�"x��S�|o���iL8/���Oۉ�r&�t�L{�)ӕS�m?a�'̃��-�𰗧�Bh2A;R���k0���:����VN��g�U��B�R�+7l����V8����x�p��lf�h?�o�Xv}��B��M,Տ6h�$Wg�}+W�P�~��yˉ��vPK��G��[�����K��X�����Qp�����g����H�޵�#��a+gF�����X��jݙ�C8���ӒZ%Ͷ��;/���U�j6��9$Y�4،<xv��;S�0}�iW7Z�A�𓄈���?�KZ���7����kң��B6���z ��$S�xE�U!�3��w�8����<»l�	{��5g~���[%�����ؠt�e��G�b��&Y�+�Q	/6q���66�7v^-m��V�ӿp����n�x$��ѕ0�ל*�HT���g>�I`J$E�����un�x\�n�BK����cޮ��PH�����Z�f�v�.���=�UP��'bA�48p;?�I<5�-Nт�ͷ���j��������$kg�?�Yo
�yn�W8�g�l<�#�k�K]
jrn�)�����������bq,X*,D���ZYi���Pz�4(6��]��I
����b.���{Q���E�*��]�����+��{�/4ǡ,��>'+6)�N�S6�y,�}a܎8�v��b������ /{�8�p��$4��w�*�g�i�]�f!u�d=qi��on��wMI垝�"9���$�~vg��[�G�m3�k�#�$H��]�=>O�T�^���8r��j�T�&z�zϫa�cz��:�ƚжݧ0�9�!E�VǢ�"�Pwا�_%�KI�#���X�ٿ����r4��hߑp��5|�3(s�N�����e���[��+��dL�:�3�\�?E�����	,�J�D�Ӡ@�QK�x����WH�^x�6jإj����G�v�����E�b8N�OX�3�(�q��2��D�K_��pvRjE�d�jQ{_T�74�E�k?|�ΒG ��7��ݵ����DG��I���H�S>�+0��R$�D�����d��gg�j�ƊUh�S1��<�z +�&�����D�=�֢0�_������o��U?ܚ�D�S-���L����d�` >���/�Y�abM��p���C��c������x*}#B�~���Ձ'���\�+(t����5��������P�S#���3��(��
j�Z�D�9V������ޑx)s8m�������
�������`�7�Ӣ:�b�۲�[��{#[�i߮,i�iʬ�^_�%Я7�3 ��!��B��UoYU3�*���,�y;�Ǉ���k?��~~����{r����	��w;K�vC�����fp��Ș��E�¥�$X��)h>vb����A��E�l�ES0E�7X��˹�O#�D�����I_zH�I�7�R��MS�y����yv����B��v4-0"IZ�5{���4z��2>DN�ϯ��O�z�f�G�~�=�:>�:�F{�^}|D�sr��w�#W��)n0��Z1�E�}��@L&��4nc^7����y�<�Ȧ{��B� !�(F��H���Z��"�K�9��.7ݽx4Sg��\�`N�ϵ ������ՄƁ~g���C/��WS �X�_+ڶ���%&��ү,t�7��p��%� ��Z
�ri�~�|B*"��rP�Rq��R4j#�1f{w��W��J��~5f]C��k��r.~�3��2��z�Z��?����3�3�m�.��Ȱ���C����,T�o�#y�2��@��Iʺ�,����j�Ӡ�g(*��l�D&/<F���H�e����|(��3�;�{�gY����]���n����{v�T��~��k��հ�!�!��t�(3vA�;�>��H�s�=�q�2��a��Ej%�j�ޞ/ J�����{H�5q�r����;��X����d^�霷?�e�}	T��x펬LtZ+%�i#���0�D+ekN�e!/���EL�n��,^���4H�'�J������F�����M`��yw�Κh)tG4p����(+#*��E��J����E֭*��b"m�Fѹ����h�JzI���	4mԝ����� �>>�t��i�T�&��*��KbS`�r~����v��p�⅟kv�Y$�m��#�m�ݟlm������9{~�����R�����1ϻ�;-�̓�	�ͻ��F�,_�K��_��;�fm_�.�f�|?0���T����(/'�d��|��3� �~/,�k^���	K�����}\`~ZS\�Z�~���K�iu�~�ӏ)�%#}س�` c��@*�0�K۳�5Y��2�Kj��0th������$QV+uUuW�ũ6��)���1�r�}·~�뇤�/z�'�c�	s/~wȔ�*!@6���C��n5���O3���y�8�ծy�ó���X^^nL�
HqV�b�F@��x�jKK�!s	��'�������g�����6q3����O�|�/�d�G�ttt���(���ٍMf�&0ڣj5�j��d��ϹvO�{�i�C����Med,e���©II��Un�=���]2���nԽ�p��l��g�/Y17IF&��IePx�g QW&�;�����'�a� K�>�F/g���@��~<�Ho�?l f���G|+�$66��U�G�Z��
�9�e/�vo�ud�61�_W�<�ݭ]Q�눿PTzz��B�F��IH��P�r�Su�����t��?�F�Ww�t�U0��SB��tl�gW��+�IC���qE˹�LX5@R��A!j��{B�"ڥ{�n!$��%~Y�F!$�~��x���-mp9w��s����8��@;pQB���|S<����G&��e��avE�;�iJ�gĺ`�H��W�۳�r��ץ���I��}���ˏ	�i�� v��`YX�B_�4,���,Vg	7	W'kMp��#`�<|wiip+'ArX`_eD�ش�W�vM)G�+;J0O�}�.�`��|vDr�U6�����(Fmf�ͩi@��#�vK5{��*n܀ԑQB�L�pwo,�E��1G�f,9�[�}���)�M��4oɿ�.��O��s�w�C��K�ل�"��f��$&�s�{��*L�e.:�𘅼��7u���BS����U�Z�8x�4�Bmv�0��;ڀ���#�6�����ￆf/���7� �x�[  �t-o@�cq���U�q�d�8��]���< @u����k��n�$�_ Üs�Û��r�������+攝_���eb�k"�/�MP_.��]#������H匓��S2�����}I[[�{������T���`/��H+0ᵅ���;�S�E&;�J�5��U!�9%A3lh Z����:-&1[�T����[hH�ܜ(��^� ���y3d'ʔY���N��=�	B%n��(��!�Z9��t�m��j�$|)�/�L�7�B��źz����=%W$$����2�@�>�M$�Rd���Y$�rJu�x堖��+#�49��Fj�z��y�l��= X)���^��"���OY��%�SpBm^�o�j�������+�е��\^���E���t��W�8�fu%��=�Ԉ��S�l��l�Ŏu��2�K�%�	<y�|��I���?�q���RVh�Ӻ�+��w��2�dHh��E������\*I���S�ܒ��C�ڞv`K��t�H�H��A�E+�Zos��������S�<[����nW��t��Zp� �z}���}Q,�(ϗ ֩ۄ���(�3R�_�eOn�4�?�TQ愠�_N"x�L�Hu��J9��YH*ć}S�dp�����3�O6� ��`�p�h`p]BjY�P���t�O��xI��I��'����y���]��E�:��VNo7�2�%=qu���.��B������	a(��W�#�̊��@�Q�����(�e9ۡ�yQ��h'�@�\�`ޝ����s&ƚ�@��W7t�!��ק�r�A���]�%�nPJ���S���hK4���1�/��y3X��,�I[����Vcq�mq�Qc�ת���NVv����J�S�~�-��H���T�a�A�a�^��j̜D��Gb�\�+�����%3Ͷ˫�y����RfN�:7��#֤��9'���x���ɣ]������̸�|OiCO�,�y�h7Ck����#s��sr�$K�]~�:�_��~}��� �Rvf���g������i��l����v׹��Z�Oq��+�v޾OW%Ѽ�z���W���wL��a9�Zws�Y��W�����K���f���#Q��#��+o> c�S��)r�ۮN��pb��h&It��$���ؿ"��=:jkBK�K\�[g��z��^�&�mP�K�H�sB�d&v�<��m�v8��t(@���'S�8���L ���:��*���H�Tڒ��+-�9qp�͹�V��$=Z�I�,��|�<���t Q���p�_��J���ěK�6B� �EE�>�lki�#��kfp�V?������ߴ�)��_��u�s|*!�uj p�#���/��B�	�g��)��n�P��ig�3������������R��@'A�FGt,�@T�@Wi�	D�\�E8���hF|���x�������g�s
��F�s��ue�j�.�5ִ֞��܃��&�V����/ �J_��6�)⟬��\}G�?���8k�!���)O�@��[W�RJH����m`E����ޠL�ߊ-��	��uR�ɜ�¢����3��ka�\NB�ݿ9�ɞv[�!�D� �{�R��ǻ>�5Q�.��s���|����!�<��;�_�#��l�9���� x�	��zmd�ڨ�ċ��+|(��c�)�12��"ӗ ���%���uL4.�9@�@�>�=�O��M;�d��V�zz��k��z6��=��"���Sj�O�����Y���c;�	��J�R���OLpМȈ�- �o����5��=xo���cN�2��{��"�ӱ�p�ٚ����|y��7u��w�){S�SHvx�L�<����4I�h��)����U'�ojH�kd�?*�Y}�� �h�i�ƿ�{g�ÅM<���;�=�8� 5�!^��}�a�$L����': �%�&�S����f�u���9��C�9G/r��{H	S��^���쑩+M���Ja�/�^�yr��nOXܫ�4\�H\��ϯ�Yð�)�<���L��O��<�~���!��?�h��^D�zs����N���kt�}�9,O�";�dL��2�#jt�܋�;jXd�a!�|����sCD���M�*A��N�}�|�`���_/�"a�»�e�0����v�Bc��Tc����M$�g������WA2�ą��/�q	��)L]�P�p�J)
�e�y�^�g�^�?����ZY�f�,��i��������܆��zٳe%��������_�� �M�;)O�a��1G<�f��>I"� Eל܂��ã�g��Y�j/�S�wW�u�7�t�H����ιlT�-n8J)�?|]��}T�}/�ѥҸ�Fä��¸a"�0�˶)��9rɹ-����<>�~)�3�K��礑T\S�+�����]��"�(v�P��^#iJ"�$"30GK~2k;�5]&	����*Yu���^F�����d^T���|��H�ۧV��=oO��Q��XI`)�k:��V�G����Y6�.�Pe`�Zd�ZId�ꘅI���U���8�_RR�1"�;N����!��b�nI�{��x�=�L��������0{ִ�ɧ'=�������2V�,���?,]��0����\9�Fam��q�?ZfnP��c��CT�qY�5Zߤ=}�7�q\?n<��A/=+2��x԰^ �������}b�Lf�U���*�Bv�L);�Z�Y�5�ji�p;^�	,��N������(��C"��z9�B%z�mu���,,��\���q�>�3WqU��2�������j~2�YLQO�n�L�̆����"J����J�\6�AB85Mq:σ6Mc�J��+˜w������5��TU��،����!�������m���gfh��[D5��@N�~�1�#�ןD��o���Dw!Bs%d�s,a+�����h��@	��Eœ(���r�R�7�>�T���#��:�A*t��fr�Q�*��ścFUa�͹��)��vm���!f��̥=�ʽ�Yy�
"��\'`��NI";��~�e����v�c�0���#���Пw�~����8��,- /u�$]����؈�&�I)N�1�̪vЭ�U\ Qҗ3�(=�hկ��(d�t	���o�S5�z)�r���R�R"D=[�ۭ˽�^���3�4	I4�MÔ��y����W'���^.hfg��;���s�����k�y;�z�b�/<���'_�
 X$��wL��\d�W�y� ܤ�C�A<�^�Ɵ�s�]U�@�N/��s��5&�D���Q�J�Ә�.ȑ��:{^~������F� DeM��n-�9���r�����o%`����Y��I�9�w�|��5-�$�**�E�4?U��ib-B�����o2��-�e���<8��z�� ���7���d���K���&�Ԃ'c��b�bF�A�jA�\�M���5j�q�1=��K阨F/S��y֎Sh٠Ҫ���xǨ��Ev���f��r#���&"������i�YQD����o��W4����L��,�#�(�־)|���&!yR��9�z��x��n���co��Q��sEc�I����Nc��8N3�������)����j�n���R��8WcE��#\s����b̬}�e�b��v�Nz�.V�91m�� �qֻ�r�����WZ�<?ڲ+.��E�FbC���Q��JC���۫/�V?>+�����z���ʶ�&1���nfNm_֜����-�԰�sLm�M�SL녚�if8�vFUŵ���k�k~{*�b֖���E����� LJ.Nz*0Pf\^&�����t��ɖ�;=�M���Դc�'�8����5���YF��f�~s[���O����;'�7�53fǌD���zy��=I��ζ(��F�e�Ȏ�=��w�E_1��K���l�>`3�c��'?���1�ǯ��(�ְu6��A#��K�o'�f0aP�3�� ���f곁����0mH}h|{S��A��ݒ�[�9/�����P��G�Pr�����+�/O�o���E�{�!D��������q�
�~-M��s]p��c�N��_��9��8�������g�^-��}3��;X��˷[!
�7_nEas����]d_cs�8�-[�Q/׬����i�
�Pފ
~�,�Ҧ��iD4�4C/b�O~��R����L���I�^���e85���|�QCm���k�������,�k��J���]@.Cx6� ��72��Wrɽi���=4�m�������37�r\��4��dlf*4f�i_$�F0��VO��N��pY�m�F��H���e��*�)&�E���ٗ/��o,G�M9�T(|��YR/�5��O.J�eg�Qy��=��`�"�L*��v�[��WW�F��)}�����#��tJ��.�5f���"����	����K^�)�ń�Y�e�E[����a�vJ�4_���~]�h����"�>ן�sJ�X���.�^����s~&�b%�;
6�I c��<������%�nS.u&@�e�z����P���p�H*�45(�'���=��KґU/oU���}+ KʮpF�7�����Y����.rܦ�%�E���gL?#(Z��7�����=�6w����ȝ�\y�3D���7�~)��9z�6�^���S�Y��ձ*0#x��.w���F������Nl6�w��|�����Gis���3K��$���J�W��us�x!��L����F�f��,WGz�J{3�?�������?��6�D�%�� ��v�n��	��d,�X�~5L��Tvz=5��t7�����TE��nm/�x�vc���y��l����5?���:=b�F״��5�X*R�k�9q:\�]j�q�U���5]����T-�&<�r��ާ�!�4.IH 3|Q���\�.���]�]�#��Lc����� '����\ը�3#\�����^�P���&ڭ(A��5�/�I��jz���w{ZI�u��ȉw��I��5j�W�l��^���3 �ȑ3ӈx��:g����G���&����/�وE��D��: �:�R��M�e�FR�_�Q�7��\�����zp�H9��C�ҥ�I(-y��kg��Y3�C$�de���IL���'�C�� Z�_�N��&���XH�s�D��xD��z���a�$;��Y��������ҽ�5���䏻�Q�l��PhZͷ�iu�����Rì϶i �|�NW�T"1>����ƾS��%�#j+�Qkd��U�`�ข��t�۪��('�W����̰Im�ġ�`�U��J-��D>�l��%+��O��8zE��u����E���`l#�>�6W����fTȣ'���ʔ=�N�'Չ�� Sm�sf��]t��b��\a����T�#�2�{��Ib��)D�JZRȚh*�z�a7�BWf�x	��
+�z���r�}�A�gN��)zѺ��f�ڴ�`�FD�?V��[�\�a8\���g(��yS��--�h��26rr�������(��������Ym�ѳ*e�dv��h[��I{ɨ������\	/rŸ�z��u��'^��t���J��4,ٿx��5W�6A�:��&�*�`�[Q��4%��ڿD״{�[MT���"t�,�*�+b���A��jWP�ӕ5�!��>�H�J{�~
S�h�3Y�.F�$5T�57ؿ�gD�˭��F�5���Z�tu̎�=��$���j��E�CL�N���ᘰt��.�F0�f�g�5��>f�c���Z2;��*г�Xu�\��o[�7�q�Q�6c�œ.����K�]��_�]
�;6�Y��,j�ڕ�]���=�@��6z� �v��k�x�����3�o��nV���e�k�w�l�B�N�F(`��Ŕ�j55%̗L��<ཹ#�ͥ��H"���;ﲬ79ӯn#�J��4<g����ɰ�,�z&ŝ�-���U����Tz�&���3�x~ś�����)z�_�HC�5W����OEO�^*�z���X>��*%���Uva!⺿$��2�b )���"l0�e%��̻���7c�F�/���:{y��O��gE��>�|"��6-��L:)=��뻁^Wv�{���%+�o_���{���!5mb��h��l��bK�9��	3|�el�ky�Z��b�$BV2o	�[y��jD�(��ѻME���W?���k������˻ޛQ���D�FŠj�߱��w�/�w�0)��i�gP����=	�tK�iιH[�M$�JP%6�a����|�K�sK�\�A������H��AԬ�V�ط��O� �-?;���R��5b�ܣ�/(����T6�)ϟ�=Ғ'j�*�s��zM-�*\�?�-:�k[�{��j������3>����4X�^q5�7z��:�l���T+��3����d2\��5�B&�jW[|�Kz+\{smez�2��$��X7��KZ(�����/v[���h��l��q-��k����}�E��������`f�`N��A����\�ppWRe+HM"AC�΋e"��@Frv7w����n��f�?E��Md��3�^��^|�n��:��=���=�]�2J\Z�P2���~q ����Y�׽T�sƪD�f�!����HR�D�URۋ3BZM�4�u��c�mJ��������r.�34�)���[R�~���(ql�2 \�jGӬ�85������;kV�Fg�wJ�߷��G�f��:��^YU����i��k��tB��5֨%`ֺ(N�?�.߶v��/���-;��rev=�jp�ތK}<5�×7Q�8(%�um���[1��=�E�1E��O��_β�,~�?�!(��
��O��eS����^V}��l�-Ϥ���Q\�+&���tGj~�xn�g�� o��̟�ǓsGL�ڰ�0m���_t�&�K���,��A�gxw����N��+V�/fVx����Un�ēY��-[tDzv=�{ Y�W��}��Fbɯ-�5��I��<ǧ�"����e�����R����7�?��7�{c�E#��K�$���D�{˷�G>2�6�C�*�ij�p�-�]��Xad�C��c�?$QGY�(s<�����ˈO�'�d���X����q�U�����S|D�����8�mI:cQY��̼�BM��ب��o�g_Ҭ����-}pۛ�+���|p���*37�.�:�Ƈ���$8ު8�B��X��9�>���|�t�#*�s'�m���ճ%�Y�lr�� Ɯ��3{C�O���֩F������6�4hح{\uHW5�=R�i�����m���g%m$��~�R��s���C���~Q���
�4��n�R�G����L�	*_�."N�M-��V�s����p�U�	��;�b�J�xp
�ZUe�j�}f�/wN?��5���#+�:j�rx~�=��YU��_:$Y�)�8��*�£�@X�����1I�*>���<�w[-�jn&N|a�s�I?M�_��Y/�d�j��3SX64u�����!�燜}eM���^�U��qB&���8�x��V�����3,�Դ͉�M	b���%���xGe���^��ON�MiZͭkb�$�q4�\yFs
��N/�du��� �
8��M�L�q8�X�����zH��3���R��z��e7M�Q��3�Zj����׍���Q�@Rb#���~��ٓ��[[�OZE�³��}OϞ���G.D��kZ�<(���"ݐ,f���4 ��b3I��Em��x��2��I�D��U?m��Y<����x�nizp����*��ob6'h�'��^��I�I寊�i��=�qXX�ĠA;�U�e�\6HL�+������--ĥh��gL�^P§�fc$�S�6V!��?���(�<T���OYz	��Ϡ���t ��j,�����	]����y�)�3T���f��dJ�Ta��vH��GQK��Jn]��FL���".��(�;���׃�y��j���n4Fh�]�_Ӳ�����x����Z�ɪ�^�rv�����`:;v�q�||���˲�H�ll�<��Hnï��]7���͚9_٫P_�89���yZc��M��gԡ�l�>����B��:I��݉�'f�7W{��M��bʿ�L�ge4�G`O+߿�q�Q �����r����/o��"_p�"�&���&�4�S�>k�*��ϔ��MC���5�N0	��Y��Ь[����O�3J,�K6�n��;�������5��DT ������=S��d���p�B�Q�c�S�_��G�ElA�|���b'��e���M���'5zΉ	�&M���ZG�IG����,�ɟ����Z�G"�b~���w�)�,XO���5p���X`�%7�R����+'��VY�P��%���cSCַ'Z�8�l�;�g���!�5.�Va���Qm��<Y��<��،>C��}vA��CC{x��*� �e�� l����������Z�ʆ�	fW��(��}jEE�ZT\;GN���ݻl�
��맷� ��G�����,F1��`V��
s3�� ����s&�F��^<W��&S�$M�dw�?y����������oZ�5��n� H<�L�����G-�l�<�zU��N�ȟϝ�}�ܿ
N�h�8��� �#�K(�^�����N��Ls��D#������8���iN4�$n8E#���R���Y��Uř���U_�4�q>��_ZJ��H�r��J��i圭��iD�S͑�5FJ/֩�+%�D�O�d{�{Nώi�9&E�F�E��Rc�xn�
;1cc�	�m�i<,ad?�h@�	��r���S���Q�}��ȟ�;�����X���3/]�RVFƲ�&��^�gŶ�iw&��0ă�G�-��z��Yۭ���\�SqW�{�߄����G��L�j-�l���UL���>���N�%X\��`��;ZyF��ŌV�:�y���q��pW�?�x��u��h��`��Q.�?�����	r�`{D�^vf����*�E�Y�k7��#�!��.kˀp{����ʧL�~m���,$����ZW$�9�h(�>&N��;��6^U%٣�N���%���-�~�u�Y���$�=���� ��"�����`�'�G�C���>���f.
S��N�x��$b�(�޵�ļ��fMڣ}C�=9}:�v,�O�����ƃGO���̠�)�#�ç�f+J*�b��F�"uJԮ_	}��nj�uV#���]%�.E���@�53X�9�Z�xi����n�@�ѱ[���Qc76��9��*�@��*]\�'84�r`�K��Ց]v�~�lA|ư�־˜Ub�
E(ILnN�_s�����Ƣ����Pm��D5h�E��ޮ�V��i���M�Y���jɇ�zi�<X�w���f?����z����vc�anf�^< h6��ϰ|_�V��3�k�r�(Y�ҋ�J W��?���Eg�O���(a��
dH�#_S��
fý�"ECbHՁN�:��AVL��L#�v��p�Xw�t���֚̊b+ܣ=�31�\�����KϮ�M"�|'�h�g����Ivw�0qԩ%��G}(Z�6#�:��-�q��y0�0��O��_���{~�_��F5�6� �m�^��+Z����3\��lO�� ^��g�t�\��j�dİ��b{�N� �QB&Q�ܿ�I��lS�IP��y��	���^G�����k��D�=v]o�-�c��G[L�ݨ�A����Eb�Sv��؜�GE6���½�����y�;;g;� 4�wE�z�Xy-1-�Eu4�~(�Q��`zl�'-�
X���4��`+�)����<�+�H&�i��4�x�����Q���d^���va�Ƣ^���5ܨq��H#O�)��������#�uPb�xH}h��"g�w��H��Ѡx+�)m�� ��y���5$�l���?~y���frdDo���2^Ջ*3D�S�0 �k0����KK�'? {��Ta���"�Ǻ�"��8��ou�h�!X���+P��O@���&�[�}�;{_S\lD�l>:_��
�3>Ϳ�|r��"�8�le�1{j#0I� �4�k���M�����v ��º,�.�9j���նf;5�`���d�l �2��w����K��mYO������/T>�!�"#���Z�����I
���O^?R��;Rq	��z���mr���7[�ۀ%��?��ߺ�0�V�b��9��6�J#��pZv6�G?����C�`�3ZrPAٻ��I��$Z�#M"<w�-��f(]�����C��0!z�n^�Y��gg�Tc�h�#��E'�������Bn#���I���x4^�(��Nڻ�z[�h��^C�Wo�$X
�����T�}Yv���*t]ݽM����_J��.9*����������eVf�2NY �/<���p�}׷j9��3CӐ�N��9�ɻ�,�0����iX���O�F�ڿ����)��>팆�~f_ 	dSn�:ܪd`vXf�x�%�\!�>�B"�0�����A�R����;1�H�Q�k���cTORB�z��̷L��^nv�ަx>��5'�0u�Ā��lBW�,�
����<�m&�:Q�`��M��g��u힧L:5X=v���ƯN���a���lA���x�w@ߞ�9��:��A�"	��r�X�S�Y1ZaU��zq+4��6(��݋������fA�\�3�Y��.�ftl4��MGpQ>��>h��:�ԘV�k_���׾��C���ON��)�hEʚ]�e���e0�!���,-�P��c��+2�c����c섌e��۩��\����s]���]�羟�r��L&`NZa,���6�յ�?��N���b�����8B{�����(�}�����N�E��uog]�Vd�����%��>ĭwBw_�G���އ��UT��h�Wu���M��D�1��Mj�V���Oy��sێ�3���,�^e33�l�IT��I�|�����/<Q�N}\FOr^ttc�&�������w�Un�G%�%M�m���ѧO����+1�O��"�w񽮮�K���a��U-�+�k�����$�Z.�tT���+�ZAs�`���G1��l9KӰ�hc�W����*���>��b{��2Bi�4|��!�]�"�°���f���Õ��Ϗ��j�wP���e}㏞�P���l~���Ş�#NFM��|�zLٙ=p�Y!]��k'K���ɓ;�[��N�1{u��-������ez�ͷ���\�B�ڍw���P�>	:���n&�$�e���ЖRr�=�A� ]��?�8@+��nc�)E �{F�6�z�8�s��G7�jFt���6>�>�ؓL1Kϒ���:�aq$��������u4��e}3g����Hr�sk
H,mV��!�8)Z:���������,G�/�(Nޫ�44�3����A_�>X�o��}�����?��?{��Y��K�����Ԁ/>�rq2�@�X��s��L*�NK�)Ա{�h�^��1A�_�Aίu��+Eߝ��ɨ$�6��}��JJ�	C}�)�lS��NGEv�=٭������Ab�����H��������9Z�W���h�׮�w��S�ڟ ���RJ�5�/s��k���a�~�s�qYD@��E~���&�F���9�ۋ�-qZ��������//o4���<�ZtQ&'u�Äg{�!�lo��&X�)�LC��JR�t�;��Kn�˫���|7\�
.�`��KU����U�6
N��)���S�H<��49�*��e!�L0�_������z̾6|p�;�
S��=��I_�.���?~�]a4Nܸ(��Q�1zS=�WW���C'��"C�eS�c�F��x���m�Ff7�G�=ğ��4	�h��X��<w��w��E���kȋ���E�;��!�u�w�Q� `\�:چ뱇wo?���UY�P:�jZ`BY���O��qv�Ô�<z�#6�hY�
�ש�D�E�{�΅�0�'��ݴ�m���(��d�FT5r��+`ۿFTs�ΘY�w),r��N��tr�e`<v������@��gܯ��q�E[sJn�㈮��v���-�����=K�fcW�R��/8���^�����HE˳LLPӫ��T�F�)���
�i���%�ǈ�~J��s'�${��\�q��g�L��8�3oD��z�Z��:�Շ�o�T��"Ն�!��0�|`�x)KMIO�0��9���T1*�A?���6��hqH���s��۱�=2c��w^�t&6��⡥(�6=p����7,eufDuT5���!�F�(��������<�U�����v���&u�'���]�MC3���m��%u�-kNɌ�P���!(\=[ÅKa�����F�Y�Kg��k�J�	���.ƏE~�^�1��XS�}7�������Q6��v$Tݏ�M�#�R�����9"��G�=��3n3n����$Xd�j���j�P���/��m��Z�lы��Jǿ�|���Cg�l�z؎���?@�Է���m��y�v��\�G�[�G�}!Sz�BI�ЄL�7��#RVIԽ"�7�k�}�Y�E����f�/�?=�Շd�9��a�D�F�|T��������>��Ј�Y�5(�ittޫ�l4X���"������AO,�PVɥ��da�[^D�{,Ƣ���dW ��0��Qswxҧr3��@VYI(�gs�{T��6, ����X�ߐ��ho�	�/$���B�D�?�oįq,
k�Z�?��7��&z�E�1��۸x�*��3�wtG�����;�S�J������x�c�<[ҥ9�	�i#��<�ц�����`V�q�sU G��0�H��֖A����J�:��C�@�5����Y#Ӳ��Z,�p�-��I��;�"m���$v��2<d�7�/�>U��b{��]]ɱ������hլ�%o�����d�;��/1r���Cr��+.�Ʀ�E{��:� �9��Bw{���v��ЃR,��Z|M�6��WN��}������rk:}�z��ڼ��l����Y�������>���d��߳���5�Mj|!�@Q-P�ۡų;��5�<	-h�,K��yM8��0�@}͟� u>}�)�ME��`P���oz�-
k��:`(ix'F�߫�"""�jf��Ij"M2�B$��/��P��3�J]pC!�#���m!Mf��*g�?̍c1�\ c��!����xO�r3�.S�5��I���lRگS��.��N~F,�*��Sȷ�l�*�)��Y�l����	�L����{B��K�y��a[u=�f$�e�d�&FWt_�-�_|�X��8~Su)ㄎ�0l���B	g�����E�.\F����� C΅9������z�b�r-�RD��o��QDΥ�E��) 8E�b�J�&��69��T��~ź����KiCN��%c1G�<�F�$�ʬ_x��+v⣗\>B��z²ө�h|��� �,ƀW����3�%B/z~����]|i#U�1��)6B6`�}/�� 5����%�j�O�11$������yC����o�9�,֣Qo�hZ��@���N-�N�Jg��q� K
��:w��}b"\�9d�R錡�+߈>�R���kg��h@�|�$g�O��8M�K#J�V<��4�o'�#"�2���KFdٵ�S����L��/�ݦ>��������c�$`N��:���`�[lC�kY����Nظ�O�XMN�D��ҫn Ɣ\ܯs��A 3|]X�髎Y��,���K�&������Α9/}�'�ɭ��ʭ�Ԏ���N�`�����_�}��^/I���ƪKm�v�l�3�k�c�!�\��s�.��KЁI3�����A��2��5��vIy�Y�_�E̫�eIy?Ϥ�l�e�:�~`���b�v��Ȧ��ɵq�� �3�Uɭ�?(f��1�;���A�u�.�Mf�����Gr� s낙��smm�-t�Q����=e��S�%c�k�3���{.���������/{��=fLm��+�~1��9�2�Nc*�R�ţ��o�9� $�i,�#�rӢs����e�{��o�i��&}G�:�N;C�8�>8����G����d��c���ܿiM1-#�_I#L�&�UB��� lk���X�,t��d�D��lh	k���y]v�z�<}Ǭڛs�;CkY#\����}��gs�z=g��EM����V0�٥�Z�Kך�����.�g��x��c��^�w�q�[�*6�U]g�S�Ig���	Ȭ;C�D���?~���ml?T��9�gR���ǕX��-vQ��qU^"c4�}::��[��eɇ�D @�^���Xa�g~�
�g�����H�v�ݶ�N))���:?%��u��zdy��-QQ���`?ۻF�HC}R
=��]�����h��<*�D&wմ�U�Im�L��^'�Q!+�l���cQ���W��]�%1H�m�L�8�s�<�v��͜nk.�� ^ ��B+�-k~t*NWx�~����h��v�.�4�/a��9>UG+W��fz��F�#��˼�,�X�D��u>䜍$�o�up.��02ˠ��� ���4*�VW���k�*&M�;�_u�W��K�2j����Z�,�5Z�VKI��:��ԯ�rWCu]2h�pEs�xk�pW��4�-CyX��۴�r��`u����P�'4
Kj��I�b����`��ډ\-��U�YK+5�D�d�?'H�'�:8�.M3Jq�H���Zq�I�8�%�Ȕ��ؗ6�DӦ�W�k�Z��)c��g��Ք�$�\QΌQ|CN�cV��dZ�b�[|��sIJ;���W ���%J誌�3-��Z�Dz_3ZX�U���n4�B� ��U���`M3T�m���@��yǗ�ΰS�������¬�Ii g�30�@���9?���S�!�`}��\#J�Θ�l~U�B)A]/�3[�߿�j��bP�U0�z+���"Û��Us3��W����h9�+4�����)�*q��A�Pz�p�<p ��*$�r("������'�BѷO/�$(=����GA*�10`׸g��7�N7R���[N�V]�Z;�$277'�F	V)K&��<��_%b-���I��<�c�+qD)����~<�4h��Z/z'���/���'����C.���Q�yG�C�r��~��%)���ωP�%3i"P���!ӛ�d�����������#s�܁V�,
j��O�p��rԳ'{�q)<Ô{�rd-۾�(ֱ�y�i��H1�5
4�I�䎶X+�L*>�hue��i!^$�g���_nx�b��%:}�{��M���kO���h�0Pؘx��J4M�4���kO(n��y3�V>����=��L[]�v�j��z��H�U�Y&(�4_x��� �b�c�F�K��`Zb!�݉F&Й�l�e����|�a4��5��ajV�B�Ky]{�$ѹ����g[�Y�������x���Ӗ~�<�L��X���Zm��o�j-<��[�#;3,w�]���<�~: �v����!`,(e~�*p��R\�'��z3�>�RW7f�g+Qˋ��Q�<������6�fD�<���~\ś��%�T27�(���	.�T:A�ɞ�e*k*�Ů��Z3�TPZ����$�5�ݳ]l�gF���9~5=����V3	�ҝ�E�.� �tbR�xP�M�|��_����I��]J��r����A	�����J��Bt��^ނ��B�`j���dmm0}t��w����^A�_����q��~����sx�~w���2��q$�#�?;��� ���o�s�ƥ����H��[�/��Gp�U�x�)���H����r�>�S�4-��Nv���mE���-%�_#���5lX��~�{/������[������s�m��I��{��7�i��]�u� PK   �A�X'�Sz�  m  /   images/b4b7fff7-3733-43f9-86f3-7eaab1c92eea.png�WWP�E �$�.��(U��TAz/�J�.AzI(FRT:"A@� ����P�j�b@�����>���93;g��즚�2�x@  �Y_O�좺_���"�\� ^`��m p����ma~r�ޱ	5�E�{ P(����o��K��L@���-u �対�-��|r0�����|{22SԈm�����J0��d�]��r�2�~�:>������OT��9tW���,&Z��IB)����Me�iQﭹ/��G�����vѩ�6J	{NԜ��O��:(s$|�T��a�k�W�jjn�cX��e�!|�1��/><=�Q�����uu	Z��y˜��{����Z�xc��8ЮP!�Pݏ����]��J�x�nUz��tY�KD[N/�!�n!h�t�-�)�ZT����HXQھb���3f����cn��r��:����?L����m�?����#"�_B>������+ń�N�O�	'�a�!S̡�ɳ.?�K�+糮_�1zU.D��R��s��LM>������IZ�Uy��N�ʻZ�=^1����&��/�j�{~�B�6�$.��h�	b���K�
�Nv�5<�5U:�ش��ґ��]|dӏ`U�]g9N+`��&\g#�&0Ii�~Wi��qF��G��Z�ɻ�<��=F#P��{�q �?�(/M�fś��&����ؖ@��9�C�L�r�KV�%���gV3)"�r���9���A�1��K����&�̑~G�ZS��`����z�@������2\c�)��u���fY�U���J��������t����N§��r��n�DT�ם��I�4ca{�4�R�/g^�Z΀����*�]����6��H����4�����ђchw�n��In�9�6s�kž���s�_�q*�8lJl�$�B��J�^!���g��YGTW��{�Y�Kv@�~C��N��p������:F�I$�y/���=��}e���!7	a�y_�,D!����\~��G���1K���۽��P�1�^���K��]/��gi:)/DT��ձ�W��4�e�����׻�TP���N�Ĵ�{�|�~+� ȿ��TfT��_v�]z6\4�^�(�/�?+r�^�-�R\+�d�߮��`vͫ��I����R�2���#�:���\���/����2~�ޞ�6�OT��A+��U4 �{��V�n�L�9]	&u�Ê�ʁq�c�IW7F���&�ڿ����:�}؆��٣��C�ܚԟ[k�&��>4/irƛ#r;���?��!�:�Q�n��j��p<�@B�0�?��`tty�j��~�✫~����]�͡����}�`洴z�hw�S@'2f  ��!=�7��r�\�pW�쨏����C�����xI�����TIΨ���Q
B��������������D٘!��|�^���t/v��_��M�����-9
�ںmE�m�K�
��{�(��yw��2'�y�4)K�	�WN�4{~G�"��p�^T��W��z\O�g�Җ��N��?��g�g�a6j������o{��xq�VD���r<Q�R�.Fw�����X5�͑�wQ�d�@�ݕ�0(�!`�5�6�8�.HלI96�<��X*����AoV��W_������ɼ|����.$��ڎi���J��Σ��j?��1��Ս��tƛ�|�;N1b��3c	e�~ͭ�W3ɾ9�2	4�';+�~1?מ�\np�E���@�9���4��V	b[>tҗ�Ψ�\n�O�G���B�$�ܯ��l����bH���r�(kDJ��o��������50qu%�Q&�l��q
ah��B$@��T�>3�=�KR�a|D,�'�RD�7[w��p�e�	m�`#6�-�z��/�R��I�A�S�ݥ6������H�G������׸�<Ի�}͒A��)��?iS'۹�dq�@0�p���s�uD�EJ�~=��[����\���Ű�˺U�Q�>�N=�)ߡ��h����Q�C�t�V�g4���5".TkN�l[���?`�z �"�����9�� ;41�r�0Zv��͝�9��E����hth��kK��iea�a'v�/IT����"�R�aQ�2��Z7�M�(�@�8qf<	҉x;W�+�\l����?��߫�å��^-MW��<������:�[��(�Q���h��6@�2zP]A<,��3���F��[��~��6͂�J>
өQ�Лw��z����	8��/���M�W�n�=�ѩ鮎(�O��N���'�bSK���%��C�L��M*sޞ�嚖?Js6�.Hz#�o`�]�k��Ӑ�J�}�gA������N��[��j�
���&�u�Z���,4K�:&��V����W�����w����'dӧT(��ϏvpI�1"���ԥ�[�N�C����l^!����d��[N�\�������y7�s�������!/�B�'S筱d��(
�f�Lc�� �ϕVG�֜�y����Y�W=X���C=O�x�?�}�Ͼ�T8Ab���'�r�}����+n����o�8�n���Q�8M�ubC��S-Wׇ��Y�Y�^h��K�[���y'�>0B

�U�d��� �.Eo���v�[W���
��mYe��>=Gc�ְ�36ꍽ�J=�U1eR�ѲoR5�q�DL���>.o�ps���t��&�V$�P���s��H�3s����t���kJw�Ɠ �K��YK'}4�����N�; n������`��~�Py��S>�_}�ff���{-��h�YwaPg���UAt����#�c@A�τA�5G`��{� �'an�')�,�8��&���2�>*BaW�c�C�t�5�0m�niz���M�c��I�0+�Ԭ֢7��q��H��d;�s�~��q� ������83�{�h/�#��nC��H�߳���v��M.�����l�ýM����,{�	�!b:@��LN`�gIZ�I���]�MK��͚o�/ܨu?�Sj��Wbo�	���ԠJ�1/f�S|����ۆ����VL�
��d'�ߩ�y��
��:n�P&)����fb ����T��>�W�Ŋp�/��>��R긥��O�9���W�J�W;�Nff��^8%�Ƿ��R%Ґ��&�YBi��3����a�����r{t?�)��⺜�D>��avN9��/:G�
]���i�alMzy唣���>2=v��"�DD����MG8�IYfڑ@:��?X�:��[t�<�MT��h�v#�lk�.��k��j�i79N�n-N�Չ@�ۇ��%
���!ˇ��&�M�i`,���/���;q�t�쩉�%��v���^���`5��o�½���gnΓ���W��������5������+ŗ#S�k�#�g,=(�.o��?~�8�~PdbM��z�S�Q���i�v�o�ք#���Y|�n���xSS)P��Kq�1��J0D����[Z��u`��Gmo�$}�:����8	y�;���7{�?Lg�w[��w������__��;�1A���M|��gJ$[ܣ��w��{��M��&�-VL�FB@�L������5��_/D��{9�|e��\�s�i|mx�S��9i��X�z���R��%�sہ� �1�l�]��5�^� ����ɲ�5Y9�9�M�G�V�׹�{����Yc���7i#���T�S���Ų?�D��^�ˌ{>~�!��82T�;����ਊecС��D�S���W��X��L�/PK   �A�X$7h�!  �!  /   images/c6364832-c854-438f-b38b-75bf2a0cd33f.png�!މPNG

   IHDR   d   G   ����   	pHYs  �  ��+  !�IDATx��}	�g��UYwuuU�Q}��P��ò�[�c3> ��L�L0��%v �`� &�{�e�X�;,`X0�c{| �u_�:�Շ�w�}WV����է���f��������������T,��~*,���t�4]М�k}��%��n �-ȡ(�a 5n;*�t����I��p۬�4(�-\mPh �����	+�~'�oQPNľ�i�xcx���Ώo�ƽ]�hvP�i �BQ�vBI�M�O�os[��ǣG��Z��):���H�Wj1
�&�&y�G�P����
l�]�!��kjW�v�!⒥vVjg�/9j�c.;�S��8����������Z�!��Z�r�Cn���]�(�v)��dE�c$ wQ�e]C��p:�X&��ܟb���g�ѳg���ƪ=7�vp�"Yj�͛���4��2�ES��t���#�bzj�u�PU��F�q9�ZU�h8�d*���F
����6X�ǋɉq4��L&O��pX�V������ ��)d2��7 ��c��U���r	>&@e�譼�l��Oc��;����u���F���N��?3����&\nL��C�����!��#	����MG�[�J �ӓ�SZۺpr��H�?E]��e1�Jz��4�,X����n��>�~:��~�K�"���~�z��g�P��Fs��� �ɑ����,l���CMu���MN!�&�"��bdl���̂������ëZ1�A�u445#G�G�g(�NL"TgEU��D*���I�Q���(*�T���pvzfi:�]K�P�6��F��'\��kUĉ�����������D�����4�����>�������sb�b���ghc�&�2�[��_�gn_U�	�-����/�J`�e!s5�w/��6�MiW��������9��V�}E(Ni[o5�vˎ�R$���������Ϧˊ]{��,�S���'X�@M-��ד頾��m;wR3����]]�kE8HJw�|Xu��6L�2�����9��2.zf����ց���Ј&��I W^ú���zNim��Qơ��7�$��Q�Vw��K�x�+aH�/��D�ӊF�!��׃�-f�^�����6�0�
�Ȟ�T�i��b�#��]{����ؠ>�^ ��yltR:���������TN��Ͱ�%V�l������D}b�^ ��P�!E�?I��٭"<S9�G��4��Ժ�ই��E���*8cYN:_A�K8S���������	�T�@8����Z�FLq���fY������̣�e�,�8�����+e𙭝0�a�� Ǿ���*Ih��!b���΋VX�T-���܁�;3q�ܕȸ|�OC'�W�"@��\�7����8hGM����?u��c�L���at��X�ž�!��u蟎b8G[�_��|4��σ�j�ʹ�r׭n� ��DWc�^������Xa���&���i��n�h&b��������p��)2Y��n���(��0ZCU������R�St~(G�cS|t6V#20
�|-ɲ�&��޷wv��K'�\��-���/"569/Wu��yr��ܻ6`Cc-~�IK�tQ����a�������Q�`��8�?۹��n��p��ÉuV�omD�ߋ�Q���y1��� ��"i�A~�D��"���z�H��Ɉ氆��۸�p8���ؗ��@i!JRʖ A~������훘�1��EX&#H�r��
��9'�#�]K�3u��dV��M�B�U�d�tznT�gת:��;���_CX�;~����UȒ�fHz�^?Ԯ �������&���!	{�yZL��Ldɜ�p) K���5֒��[%3�����;G>�FDIҀM�SD��``��찘���!����vS������/s�� p�:Gj�'P�/�&�M��i7�nchb�f�@)G�Dc�Z$�ŋg����I�Tx�:X��3G��O���
4��&ȖO�T�J�w�ā�29�R�f!O���T��pD�3���H
llO��g���J����A�|��Y,��q�LG�$5AB½k	���e�>6!�E�p�(����Dd38�~�)������89|E>�%!a3�-1�+K2䏫S8�y`3����h0i�
=��*ND�񲽎.Ē%FL%��$�f0��y=�U:pa<%���'F��T����Q"3�0d`�/Αy1JQй���Re�G3��q��_��x#fHһPi��3׍��Hr/E��v��}�E�H_�}g�_��H4�
�7���^��&�7�/|�3�r:�����Q�mU�R���J7�F5|;��hO�8'.R�މ�t�U��6���cf�.�Fj=�'��
}�"CIg<���k��i��XZ8M��7�	|90_{�Y&�R��kT��X���cqS�8�`Ma���f��%F�)
�@b��͎��o&~���^��b}R)�~�����i3��[Ŗe�d�6{��2wŹ:?̜6aP�HD����Z����8�:�*�Đ� MQV�� =݃H�zd�������)�T��i���
���0m�n�m�ߪ�yE��ܰ��R��H����,6Al"��EÊ��!��33x���}g�Ŧ�}�!>����^��߿��`������f�q��9��@w���lz7]#g5s�����M&*�)�e13H*�>BG���)��ό\Y����m铲�L�M|�Z67L���c�3��i3���%0[��^[W����3����;���T����.m،qnB�1J݂����&Sf���.�A�b��� �HI��?,�q<�f�M��#�j���6F��$�	_�4�N���_&ЅXɳ%�d�&����KOh6�ia�3OJ>�$if|G<�t�%y�|�d��2��Y%fVy\r�	X�r�(0�����'�e�)K�+��Vg1��o��;RrZW��2ODy�3�¸!��
��Y��̌:��a
(�9�ϻף"�	��_<�,�;O�.�:,�;���={$�LPd��g��[��_O���ޛqφ�T����'��S�"���6Y�_�f�:��x�#V���9��
�6��O��i�_�TpqYy�J��gfwi)ib�T�n7��8�**)y�![�#����(��9�է��k����������ַ�k��6������|O~�����>�<N�Na1��o�h����I�vܷ�/�_ ).P�8�5uAѲ�(9�g�͉a���7v� �Ç����s��5A�����z{°��
�;N�G�+n��+2�W�,�y[�����6&��{_L�*k��g�p����?�߱A�;���Dߵ�_y�5��F�v9(b�r����V�{w�7�w<�OߺYL3�����%ʸ�.'��Ղ��g��˓��f(�v�QM�S�mg�r�;�S✍33Ù��y�1�Ḛ��������a>��w��|��Ib���~���q�??&����;�Dy�NSҹ}U�� 9?!�R����&�Vv�ϝ�~����!��5�)'%��p�n1W�f9�˄t���;���g��`&��.:XӾ�g�,��O`)e��&��9$-w�5b߹Q|���bj�8އJr�~:"�񼝋r	6�����lN��a|����>1�E�*���}��"�eq+O�q��eO�����T�t��4���@�L&�a''j��LL�w_;���s�H�ӽ�"�~/~��$0����>x�����ɡ�����o���i
8*ȇ���,��5�w��sz<�f�O�~6i��L~���)�oG�bKkz��1�|�Qr��n��l
�N;O_5��={:����	3"Q�kM67Ւs�P���ϒ�'v���i�E������I]f[9�������XC��~�%{��Ħ���������\�W�>�g��)\Of��������L���������DX�88`����Z��x��1ay"��hR��I��>�έ���-��()��ǑD@�ߤ)bc�V0�8�i:6ӱ���WOCs:��o��M�����H�9�KĲ���K�$>zC'�m�R�x� ��et�cPR�D؟���Na+K��<�~r��0�CZ��_�S=��]2M��C�(2�EI�����'�%�[]���5V��7J�������sp��Ϯ��m��ZC���FN�tƇ��G�Ã��g���׷��J������ꁫj����aUE[f�(7����Ȕ��(U��}�~�L�a���������x����)�1~��*]v�b6L�C��?8.����&�;ֵ���\6��'��j�y��(�0�Q���B�"_��,}���1�e��O�|����{���� �0-d�9�� �:�Y���DZ�ſ�;�H�\�����0�P���3�s��}�u;�r�whxS�Y�3s֞����	?�
�g1����3�f�,�2b3��9;�����\�(���KG9�\�)/�R�"�&���v�!��N&kϝ<�#S� x�-�cUx��,����|t��qe$͉K&
;y�����7��P�1TY����_��?�c'��O�V�U-�G�lUf�후1f��7�/;DժcY``���RT	c=�kJ77����?8���LV�M�Uʢ9lu�VL��U��*��('v���+��1c���1<�8@��a��t��m�5E��*j�+K3Ư/�����W�%��"�q��hּ^
{�뛜i_{��sU�R�S�g����ǥ�i�J(����� �,/e��V�S�����!�ݨ�o�
��Sc���4��{&�%�%�뫊�j�Y_�7`��0���~�"�.6X`
f�,�]�av���	��<��N�a)de��%�	]
l�U�N�4-U6Y�W�MNY(a{z�a4��OMƳM�e��_z@es��@!��@&P�8C���IWxkjq����_B�߉���D�u�^$�9�ۄp�*���s�h���ܗ�?0rA����ZWZ�H�"��3SQس)xm�+01�&�VDc�#�t��W)KGY�?Ȝ� ����(��0���ݕ�ȫ�u�|�~�"r��j6`K3Ģ(ט�� I�j�n����d��J>�`��n �B�������A��	ԫY���	/�>�E��7�`x`��Q�<U��VC��g��C�Hd4:~�\�Gjs�g^M�� ��5�����"'�[�y+G+�/P��J�!�xE�q�D���6 3%O�F�3�XW��32;���Sqb�&�W_c��<�hXuEJY,<����y�r�!o5pt��44��x�@�����]A���q�D<x�d�-`���ባg�/R�ѵʂ�>���C�ష��`������5��Mp�s�o�!�L'���(-��5X�)���~����S��*��?g��BqW �鋬����+b�;�w
�fL��czP��a�e(�p�4����h/Nf���K޲�w0���^��p��&��(��U�A�r�HF���D�S��	�v�9s��J3��wbP���cE�y�v��>�f��%*�	��"2bN��L�����hЋyٵ�!&8�S�nyg�$l�y�X�2s��_��*�*Ic�;��O5;PW�ď�
x9\���+�_^�E�3�ك�D߯|DKn��etD�:��j��~��3d�eAe���ɂT��J
�5�,��f�t^�7�sd9�ȥy���J٨��&;Bd�/`_�L�5�\6,�!���"��)��y�3)r\�A	(��ȼe9Hi���Ey�-�>D_��Wd�d�P�@�e╡�RIC��{.e�M֬�l�nW޲n�ˇ�����H(9����iooG?�<�_�#�5+%0ʢ�H��:��t�>��I(���//�'"&��TS����������*?.'�V-Hk���x}'5���y�T/k.]����֟;�h�.?R���^�9ӊ��ͱ�#��=pU+nڸN
�x���8���K���P)����E[[vw�¾�!�9݇�@��a�;�)���f�[,ڮw�z��
`U�Q��-�y��RE���̓�u����&pv?~����GQ][+�b��Ə~�#|㕽��l�06��g>�lٶ�͎O��G��K�����68�,���,ʐ�7"�H�)�סZ'��Hj^ۥ���V͙wfu��ަ
����B�q �PY]�O�٧����'�R��/��ؼ}�T��
1eˮ�x��
���p*PK���wf�)â9r�:::f�s8�L��D�Uu.*�#.2)���ҥ:�������e[��~���}����m؄M7�(eYg�#�͠���ݲ'��&C}���[,�� ��t%�K��`)��w�L;lW&_&��/$/�yn����aF3f3���5d��;;.Q+DGWW��=s��L+��1d����rŋ[0�0�b_	��)
-�z�p��5���bb��9߹�z���D
(3,�~������|��\�@�bL����R�*�%�xAx�	��}���r�̮�S���^8;,E�̂2����|ny�|(��]��(�Y�
����}��$:M������*:�8ݾ�-���a���Lb�G�Q9|���=s(���NI���G҈ݶ�c!Q3�4^�u./){x[3�Ul������q���9���2Q���Uu�g�9��p�����0���C��Ɍ�]���0Sjp,���r�j��H�pr�gNJ����]�]�MF�ۿ��fHYfCAY�u쟿�u|�k_C$���0JUB!��@���Y<���bt|�d��֥��v���B��ٚƛ;�LDG1���$t�E�/�]-XᔭmRN6�Ɛ�ʮ,���-.Zz�պx�i�D�P8.�)�����'�A��q�cޟ/����l���cH�"�C�_�iQ\s�vD�)�ȡONO#�����p��Ĥ�v5����O"�JK�v��6��Dcc#��uT�r~&6�&<K'K��|�Օr���XJɤ`��2�At���|�R�ᩞ��E X�yK�l�[��ZޟX,�JD.N0U� g�Lv򲉒efŽ��Ic����N��鸑��\1���7�����d\��l�_Y�x۶�KE�\Wᒍ@}���p���ۏ��fX[6H�SA���և�SIL��M� �]qU:~v�t+K��$Ō�ON�Z����i:j��睷�q;� :#'Vs��c�Ke���#�d.��ppi?.��1���
`�|L�4��?0S��vz�v�7�R���.r����?C3��&�sr�!��^u�L?.E�C���y"�b1OYj� M�ʾev$�5�%?1��q8���&�����3s��'F�?Ra��:�/�I5_)��G䊆<�,ȩ�OFxH�:k���YE�a$T�X��&d+?�`�Of1_�a���ʏW�$�� |\7���|H������h
Vs�o��B� ���H�^�ұ����z̳�2���j�*�l��A��O��X\�X��YԸR#�Ҙ���S)�x(fy�ym8
)8su���I��Ǣ\N#�b�p�5�>r~H�tr(��8~�"�t�s���#�%A�0�	25�|��'Ϝ�����Y�d�5$���z���35��p�!6̈́#L��S�BOdq�d�
u���ӲAǫ���IL�I}����ǩ˿�t!�T��l*�*��v؛:68[��31���	?A�}�D��s�B��B�{�i�m'�������B:����)\�!�N���#)U��G�@s}O��|.�Օ~1s�x�n��Nj���e�,2��}>��}7R��<�f�U�^����H}I%��x�bw ��I?��*%$ϤS訬㯠h����J&Q$f��6��u���?#�|��[�!�<dl}/�w���b!�a���zq���dR�kJYp���YImy(g!�ǎ�su%�NP8/���-[��_�9��[���If��`�#���Ν;)�Ȣ�p\w�u� SvapP"�M�6!FAƉǱm��9&�5}z|#��c���8z�� �i��_L$O;MG#��b玝b�O�<���fT�z00:�����m�d-_":ݯ�uw�!�������t��:� Y���w/�4����]	"�ljS�}�fю"����mb�y������ۥ�-�=ߴa���		�Ch�J��;�m�v����5�;I�,bf�>�ھMp�RKc��ċ�I�wn�j��֮�܅���ڶM�E��o�qԞ�����͍(^���23$)�?h~X�s�bb�?����#F�,��_.�ʸ��P�V�-E��U�|����/N��Q�C\�����W��)yk�����[�߽�9��h�@4����fJE��YDp�g�]��Sw���n�m�F����a��7!�3d�_揂q���޸~���M�I��)�G�2�_n���"S����,1��d%�³�����1� S���    IEND�B`�PK   �A�X�+�s;  z;  /   images/f3037bb0-f56a-43e4-a2ff-17056f7c669b.pngz;�ĉPNG

   IHDR   d   d   p�T   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  ;IDATx��}�dU����z�B��=��ff��a� E��~���bXu]W�[]W�.:,b �H�!ϐ����=�=�su����ι�UuU�V�ou�Ztͭ���{���p�S^i���6���-��d~���q����n�%�c)E�Q��m2i�΅��Xi2S,��'m��.�FQ���-���Tm�����b0s�;B�~����e�>'Ax���;hW��������߾Om�P�-����sC�z�C�"�"�ZȐ4]PR
��m����5�������(|��D�>u�
e�ڶi2O]�m��$��0���9@m�������+��XҰд�OP�1,�|��� ��r�:�P�����:駙9E�)�3��5Pn�H��~{����mַ_��|���O[�)�٩����~qme����
`q���eIm�ō��!-o��/@Zє��7�dڶ}�|���m�
��-��!��he��x��u��6�o��~������_�$�.Z|��/LW����yf�!������o���h}/�|s�o5$��`qQ�)^�Z�,�̲��n�V4��8Ǧ=�`���e��J4#f4���`ZNѵ�iM4�h�Ry@��Y��3XL��Ч-F�����k6���,��LW���a:U��!�����
�<�.�0�x��N詔<�Q.�f�dw@���H�t5�C?z�v�f�ॕ�g(x����sYRa��]�^��Π�)�Ѡ�fF�Y�o0��C0��+p!�h�Iv;�H�8]���՗
 ڟ��h�4#��H���A<v����A2ɫe�{��caV(�(�Qiy����X����3�W3��@X��?�EI4c��j!]�"�� ,d}�D׮[涯�xSԥ
�3�2�b.CZrbe,�2i#;}Ƞ6�d5k��x�X�F�`��h�o\i:㼹�o�K/<��4�Mc6�*�Y1�g�b�)�L��E��>y�يܺ�652�=/�P�mWHa���H� M��Z
3�3B�����h'K*Mk1\��cC(?z of���.j�X�d�X/�Y�Ҽ���n��iE���1kD�͊��u'�_Q���n8��c�n0e��ym�à]2��ߊ�T�u��=��,�~O;�;=�K�n�"V�G�VB�zR��GV��D�q�[�Y��[.-n���Y� M���1�%B��Y�R3���������Ĳ&X)��X�X)\N���8��������{~���*��X��4#��j藃B�dY֓�P�6�t�H�����f�̥��>�Į�M<�U?!���|�}˜϶ؙ��<�����6��p҂���nz(CT��>���]���߲����[�D�چD".�a�.�߇v3"�8!iU��[ݼ��4j�9����#�x귏����c�觕o,}~�1��WRʂ܈�4�m���$/Ȑ1�6�������ӏ?��J1ޱ��,�u"1":���L��qO�Ik�Ѯ�!:�PuY1��+#1T66b� �x��)�E�z��P���ebJ�p!�BMQY5�=�@_��y����s1��҃ŭ��՚-�]��}��`�Lc�4�E1�8�hV҇6{F�+aAMezN��J�Lo�$�]]���u%P3,�)�c�D&����&�������D��ٝV�J���54���[`�B��2f�V;m-k5�uz0�?.�d��8M3ᯮ��ӅvR��OΨ�l^����C�3���'�(�Hf��,�o�&�^�n�^y�;_�n5m��F<���*�d�[�8��z`��J�`_��D��;��!��VRן,s���@g��p8PQQ!��O��eg�����)Y(��;��o�.X����ΚfX��0x	����k]#�k!;w#�3�:넥PK�C�`���:�E���=S\\�?���H*�Z���Ls�K&��H�h%h]ؾ�!<���(00�L*-�|1q50	}�82� ���X�N����o~�
�;C��W��";f�A�Ě�O���P�a�>2u�R*QP�c+t{0��|r(�F����f�ʈ�g6�^3܇�ۿV[�\d)n���e������Շ�o�C~4�r��U$���i�%I�T���좉�!��:aŮ#�#��Q�%e�����E���}Q�����<�h����4GؿEE"qv�ˎ3��B �%s�%�/- �3s��lᕖ`+�f=+��i�\f����P�I�ξ6}��-v~:����-�CH�&�|���{&Q�b%�z{�EgY�:����:������m�ɫ:��x�x�w�'���]�ǡ�*�t|�܍k�����F�UR`��K<��[0����o��zW�>QgGR�����'ahC�=�ъZ����Qd"���z��ƞy	�?7	�Q2��C&6������ߠ��sz�p����.���HX�2q~>����Iv�2ы�Ƣ/�'��g��iH�;}U�V�
��t�H��)�����0r3C�0������$��̶<p)�m�o�9hi�HN0>{Y�����E��CB�i|��jH6R}'�����4A�kj�*L���V^)�(��a���O��@�k٢�$��5@'"9������D°R{=Grt �8�d��Zh�{��TYEmbЏ����*�4�3�K�ӥzV�Ok_h�� �B�A�C�n��g�gƆ�coB��Y�����j�7�L�����	�W�L�c�]O���m�.[����u��P򳏣���a)��؝�G���!����|U�y��ct��H�1$b���gP���g2��?���J�$������-����v���'�p=���^��@/��%p�{���;܏�+އT�a��䋯��Ӆ���,�u�QMe]���G����:
^�!=Ǡ���#���,�C�����X�H�UP�e�p����lM`5w�.\.�f
7N:;(�*e�I��I#�JqzR�}�t��S��B�ij�V�DM�O�����]�@�O�~S�Q�-�
_K�*�O��Y/�Eu�?�pԏ�6�c1�%��t�sa<�l)�bvH�woC�?��.+��4�.�i�ҎE�J�5��@Z���"�=��Ϡ�̷kl4�IHU.���v��t�LP^�R� �i�T����5H�hB�:!���	!XH�����-��ό�BO&��0��#6��C���T����a�R����Ӣ��	Ȓ�>Mb��!{�P��nc�)�,>3$2��i�fxኘ�0(Ғ:Ns;q��C!��yU���S�c�7����k"@3 ��4�ii3S�y�Nz�J�X��e	v�"`�;���:�B��
A0-A��;��7"��FJ��H�B%]1y�� ��Ĩ(\OO�c�G���DL��J�[�x&�M0I�F�X�'��oC���n�`�D��L���H��hZ��	�}$@D�т�1��y����|4J$#~��I%��f�"ZS��� >�>��UM����f����v�_Nm��5<��`�D�'�UX���H��~*�#�l��*����C�o<uJ!fRC��0�K�����Y���ob�F����cV��?�=�x��&��e�~��%=
3#��U^�:���ue�8�)"��9�"��b\�~9��������i����7�?D�_nw��M�L/��M��s���s��9;d�P�=�O8V-2Z�du/FN ��_/�ȱ!�0՞v��}���%Bm��ϬϨ�0�zF�N��GF7��r�i[8](�X��uE�������$�����O~�n9c7]������Ӷ#��au�浈%�L�o�Z�E�$&�7�N�Y][��HN[��� 95�W_��	��c,>�N��w�����n�yYhln�燈����k���Mm��a�/&�Y�q=�B�lFt��z�G���0�g��9�^���f��� �iaC����!۬8���9h��=p8��$@�
��h��K������o����VU��uo�R��[i)DШ��d"���
�k4{�f����@����Ց4	�z��ڲ�O�'�E@����MŨM�\�v���k�ꢬ��xt0���T�(!�p�ظ}��CH�;�g�����,����K���Yh���!�ӱ��t� �L"M%�CX�*o>�?��C�y�dt6�����ק����g����eE�>-���/������x�p$f�8����ԑ� ���Ț�!�+��	��ʜv�=Dv����N�|�KA���7�B�1)�ljNQ}�=��;d�!�H���3��=���@s$�K�feD�f�C$FL/ll��;����V�<��7#�XN2�˕v2jB�˝�@�����D��k:��߷dt=Nl�p��\�5&�tQ%{|S��3C�sP� Ms�Éd<1�������d,mY��7�wS�_�wi�w�4��~�~0������Oi�Y4L���%�00HD�&R�F;�s�"����*��;�}���e����v���'F����f�&�_}��}�:�Ēp��������n�IcwN���:�r2����l=��X�픭��２�����׊>؅�������쇢1d����1r�LzA#���(�"�P�u�[�!,���сa������rܰe�	?��r�B;�Ey��a9�t�cU�;ػހ�؎��!A#�$��meY��s�5@����2$�	bH�]2�t�1c����\=�	v�����;��=32$�}n��a��ײ��}q�"��8��
�{��@������1V��@�4'8Dk���o���",;��-ȹz�����:�A~��ާ龳�!|����v�a�/ːI٭�myF�$��bV����b��w����A1CF3Sǿ����
s�'��?%|O�Oe*?v��fq��e3����-4���F{���>���^�f�_�������2�nN&S��=��b�,1�E�����F�B��b��n�Ӥ/��a���r�v�z&^Vp2\�2�'Ơ%�0Ek���ԊL$�����Y��U�����@g�^���#�u��{��뀕���2�#ƭ,J�}Ub�����R�B�׳�a��HRȯ��"���J���$�����
C_�sti��2-9$�)��UX��k��D��vH�D�}��C�"r
e�\���F�H�����.F���_q5��
��m@��qq��K�@���&�x2g��E��h�_��I�\04W)�Vݢ��(�{(�� �~qY��y�~�5(�{ 0=��`��P���pd4��ë��ِrb�x�LJ��W�vHn��gZ���Đ�e5,En��ȁ��\�$¿���h�I�7�#nm?�e�����]t����!�~z?�'3��hVL��(+�'�'�![&�Q�����PgL�f��~��AKP�@.f�Ёي6[��\�~Y��� ��K��ٞ"�'q�z����Bv:Qt�F���?���W��l%2�\3�r*��������)l�횋��&
�b�|6��٢������I�e2��8�W�2)5�XA.dk�������0���,>�\�[�b�W�@:�l�Ӫ�8�!C�.��]P|%P#!�D0�³(�~�����
{0�QKƌQҴI_�@xYhN4�0��� �(%�BɆ�z��"Y��j\ͫ���#��+p4��:�t��u#?���V��?�A��v��(m���b���#(��5��p��'VW��?$¶��8����Dp��g!�櫰U׊	ȓ�VY%Dw��A�ܙ0� ����m�VQE�"7��ar��L�@WS�@FB�Zb$$Y�s��1A�Ǎ�l�8w޿�E37N�1	 �z�D���C��XfxXYXD�XQ��fأ��Ӌ������G&M���`	b�ٽ��	�[��i'��:Խ�dB�GM��ޤ6g	z�{�i��썶��iO�<t@(��Ѐ�<�N#������V�
���;���$���[X:�z�ɈP��(�w͜La1�Ngo#�#@���pVz�a�Y��ٵ���2�cN�هk7��F��wb����U����H��B+�1�� �1%�oG���D�o�V��.�/��s�a�0_�
�e���3�Z����d��ayE3"yi�y�V��AݎǬn4�^��[����E�"�cq?~/��2:;;c�_V���w�Ia��~<m��Q|݇�#�X>�vZ��|�k_�/cC��=�1�G�B7�T,��A��r(ⓗ�gl�ǯ�n�:&,Di#��L�W�G�n���?�{�)���"Z �a�i��amA����Ah4I���'�4��p䅃�R�(�P,L�J�*�|�g�A<V�̄��-�i),�憢-`e��f������^�+.�^"\6��g������><�������L�1�q��V=����i��W�{��N�����&Y]L���$2v��D�B����C��'�Z�] ��
;Rezv�W��-H?|nR��6!nu�%{�T8��=�뗠{Z!�H@=F��ƿ��+�<�V5��	�3*I�S<�[u��ۧ݊+;����DҒ�2�� �ǘ�@~G1�~��P�?���9Kt8S1�w���x�[��~��⋌|�drF[�ۍ�r����b�)fw	�X�f�Kb,��C���aܶE��c/l�r��c>�b����!��C�¦�{�|��HZ�yb��V��p�57N#}L+��9,��}R'��>$��ܷ�����k�M������ʍh��M��'0�ė���-���3O}�8�u�pa8�"1�����%m�`.�p=3���'oڄ"~�9h�h�ӆ�n���>M�L�q�	����$��_R!]��5lw([�>4��<#'�K���6v�JvY�hʆ��
��꩘^6��>J����U��'�)�$%Oޓ"�y�Wx`�bC�V��eZ9�2��-�W^u��\�(Y@��сM��b�E��х�9�f��!M�C����ڇ����a�V�qZ���c�A8�[HIy��@�	B�_�S^J�,C3K�Y�E+��bS eǓm/f�*$�����6��d;_l�r] y!��?!�0����g�M��9�4pk;w ��DG�+~���tE#}�o��+j��	�� �(p�%^C�=.�Sߘ<�@�Y7Ŕߡh�W�ؐ���%
B_��͹�"[�Ղ��}E4�{C|���p�Q�dВ1X\ޜ��=�(j�:�&�XYY)`��~���	/��"�2CfIr���`E� ���F��w���;9����p(�7P7N��,%���ɺ��pVT�}�K-�U�\�>��Ŝ���0;6	�{��%dx}��_b�m/�ɑc�����,8�>I�e���R#1����*w�\(++CMu�	j��̙���ƻW�p�d�$�h�����'�R(�x�ڍ� a�A�rF����ņ���`�ß�{��<�JL�~�= _x"0�
N"�ԣ�#_DQ8���/��D�\9�+#!�]�E�2��.��d���
��p8��H���c�/ Or�I[,EQ���x�C�#�#�%��=�Xk��bt�0c������5t�n�v䈱`��K0U��g&̸'��tc�3��D��|����(��:Ay$�e��хzlJ+�EO���a�H�����pCQ,S[60�i@D�0Y�G��!f��8󯺺5U����#����h����Ç�q��֬�v1��*2��xb���21&���o3�~�, ���֞��}�8�2+�زb/J<L�4<<Hv��N��*n�?X��"�,p��!UUU���LQ$=I�B]�BkɴL�k�	��-R'(��D"�λ�����+�PRչ���l�%.�,���B3���hoG�"C�|[+�o-��V�sX���&e0���{:�%��԰̜?3z�V�ɑQ\�e+"�Q2��ˮ�h_m�ˠ0[U#G��{��̲"]ŵ��7^Ƿ�������[��pS�EL���FaUk�1����ۈ��|I@� [�Ծ��ń�M���[n)@YYg�0������,1��Ċ�8ғC`��۲
�S����E:�B�Dn'��GM3�FY4.�ˍ�d���Uը��Ĭ8���	�&�U���f��b�J7?���d�󷏡`7\֮]+c�I����}xf�s(&��,�l��l�㍞�4�5��e���@g�S"��}Y�#X��0���(��*����`���;	�T��d.I��4��@� ��P��]������8����F�57>�������>E�8�����Lx���!�Z�
M�a=�H�����µRc�#u�PS4�Uh�i-z������/��T���F��~�`��b�ϋ4d`` c��|�=Z׬1|\s0�Y�q�Dx�wX-� A���7�N�I���	T�!�h&O�m��+�*��[s)uj;��Иe�p�Y%%�������8�����~�H@�0S��q>��=�^{F��`k��\B bU�z�n����@U]����
l�Q�����"�W*.���D�*u����&h��D�z���3W��4F:�	x�⢘|ԟe�n����*�X%iى�{�xz8G�*HӺ��j�n���2�/L�"�Yb���8�&�M/̈��^�S�I[�I���ҁ�"SXI��e�S3F:�}�#���	|M9M�O{��]��4S�؞K�еե��|~���9��4�	�zpa�	����:��'�Q�NzM���l������.f�[IR�$�.�����!�zc^��Z�
Ȭ��ŃH��%f�[Ҁ6��Z"^��Ļ�}�S�np�EƲL7��PL6�H&�Ԝn�̭��s��%9����"�W"�����>�n�B�m�&l�&��<Y%�c��/��ƅ$}�<76���ǡ�3��7�� �Ua�I�����~�N6��[�R��a�<�^	��):�O��}8j+B�KAM���(F�:�*m9^�n'n�����p�ھ����Ӄ&E���2�W#zp�'���ߋ��h��ۍ`�	|��# ?��ag�x��Fr'!\'G�n>�p�x��L�-
��FFFP�~-���j�oWz!�IhW0~��aTUV���6��MU��?���M�Aó����7X�В��t�3���>�I��`�-��a��j���c�h.;����a�:Y��e�Wxx?�������=d�0�a8���|�)A�އ{t'A͙��YtG��Q�i"
;;N��|@A�P&��:E�IG�<St�2��|4>��b:A�k@(�0��DC��**��r/!}�z��ć�,Q����O�O���&K}�=��1?�)��p�s������y�#�8A+㹗;e�w;Ĕ���G04�4 Y͹]�*xq��Z��>.ғ\�Z=|P�K�rx9��l�_ºj%��<���ݹ�!|E�D���"��Jp�����&{g��{��9��� w[{��}��dk:�O�'��
�A���A�P19�uB��đ+pP��JJJP[[+���ȉ�jG�E6�<��|���R���&�1*�d����OJ�.H�z�
]$�͟��̨&��!�:Ja8hL~�����;}�L~?�L��3�!��8qa�'w�Y6��#�����_Ax�F��4�������L4�e�턪&V��k��N����Alڸ�_v�ܱ�>�(���66`���@��.�9b�X}%�^?��W�QRQm�(
�$<�.!㩟�ub�h*���j�e���+���#�����\e�����E"�|�>LsJ�M�c/��.,��`I���C�xP�_�au"�X<dHB3�Kl#�"�;���՝��34�Pz9M�Ёɭ�D��Kn�-[�o����.l�$�b����[�ك�^Z���G��P�����=�z��`��M��T�JZ����N$o5:6�[O���}b_���+Ѵ��h�x�U�2����=e;��,�d�`Ög���[C��~�$I݆h �FZ�	}3y�\YfH�~��L��$N�<�#�w=�����Σ����w�p�͂<�椩�oooǦ�N��%�}��b�5]�ޯ�iSv�p=�ů�g�^{�G��}�qU�r,�4�e�d6C��T��6�uB������'D���&�E6���14�M�P�#�1��*���g����fiqĐ�-�səL�����	#���iF�S6�['tF2�p9{���c�Qݼr�V���C���x&����g�_��ݮ���\�"T3��=b�o�8˫q4���چP,�DA�a�l4�W+	\alR��#d9��������:>t@���"�Y٧zc7���jY���Qw�����8����w
Ĕ�;Q���Rz�%����V��N�(Ny��{�J�uv��!v�gl�"�w2��+?���"�/kF�nZF��>�Bg��\�ؽ�m'��ϻ�x�`�F����� j�����
�9=ة{jjs��J7-�GFe@1^8A-i�1x_��&�1-��3�5�l=KlSQL>�4<��F�����M$F,(jY�T_����G2)n�8�H��@O���#�ۀ�@|g���+ϋ�
����!nK�Y&E޸|�����>�gt����Ҟ�獻�%��J��)���g���:Z��Hϓ�i#��X��o�.i�Wu<��,������蓄�톯_2��L���[$sv�M:jz*0�\�;׵""�<>��\,E�[o�,� C=��C����aD��`�!��@"��BǏ�H�y"P7���u?�G��pM ��S�˼�e���Fq�v.Ab�cɮ.���n#��!+���6\�!�^���$&�T1ƤQ�;t�C��=C4=��+���QxRQaq�R�s���=�:'iZ���[�l�d섽�A������u(�����dMK��J2�q�1b^�9����Ȟ�#�W����Қ�:q�
�q��%��O$MM�ά��i���x� ���	z�]n��WP�U���v$����b��P �w���%w<�˗§�IZ(�+T.ݶ��v}��O��b��^MR"J�]�+क�	؊��4{ݰON�E2:v�؎�&��(�B�f�N�׹�T�[OB���H���-kB�d��\�lTo1ĥ��2MԨ��1�Mے͓���0c�o~9p� .��,�P�n$��;O822��=>�.���J�:W�3!r`/�$�#���ZS�T$*�a:[�����!��4�Oı1��/�U�\���~��.x��Ι����v�vثV������?*�Qݼ =|5�����q�kP^���ŞF5F�՗s�#���{ϫ�QG��b�J�J��-^�3���J������*D{���E��R\����)	fV<����N������b�����"$߽[����w�}~�[σ�3���?������>�?R҄�n����)���	f����[�
S,���'1�%��r��r��mr�K<��r�6�S�y���c� 4;$�8X�<��� 0&i���?Ɨ��c��|���ouu��F�ܫp��X�Q���h"�,��+���z߻Cl�)�~´J�6��!!N����9
�(Ь����8c����/�燂�V��Õ��V�E�
����bqó�\A\�j���&�����w�,2��kk���l����ϣ%�%`�d��0�����!>�����y��D'�����w���s��>���p:��M����[��Zojj��3�YGɱ�����[k)�+�ov����Q>6������4����غ��<��X���-JHS'�H����Ŝ5<uޡ.�ϲ`�D;���`ǵ�@��Ni������POn�c~"C�H�ߣ-�{xX�>��?���ċ�}%#����
��8V�g�Y��8�ÿƱ�n|���ओNY�<Ax�d0�ǟ~/��Cv�W�ܣ͒�Ęs��/}5�ӳ;�����5��[��}��nNv��F'o��ྀ̽s�y���H�Q�;=����[}����H)(���o5�!��J��H�1�ɨ�Bh���0"�Bm_%��co�����W�2
�3�g����뱬��'wubt2A"vj�q���"S�"�p������GCC�4�]�������H�h�T%��&5Ǵ�[�DL�N�\V��V��kO�ˌC�/��T��N�J.��.��|1���nCI篰�p�8�)CW���KkE�n!���`�-��Ѩ084�~���wC�"]B�L���g�j��z�2�#�ܗ)ű�w@"�u*�0���7� ����2�f��ĔS��X�j� ��{L��s-湓�D4��]9�jxz�{F0H�т$=��컛&�
p{��Đ�׈�-�rbf�<x�o�ג�'S�֪
�%xxx�ؕ~୅�>H@`�.>���"�S���Hv���a��˅b�/3؉u��u�p�}⁹�����ԥ��V��Hb�}�rk������$#AB���1O5�����n!)Kbq��xN^�Yc0_�����Z*�X���l�t��!��.���^ ����rb�˛��ݐV4s���,^���&^��o=.H�{HR�y�Z��� ���9�u�J7�у��Z�hʐ��م�"ZeV���4�d`n�Ԍ5��3b�F��S��S�� ��E*?G���P������˦��=4�Q�ԧ�:D�w������01/.[�=0:�	������II�e����i!>�ה���5��$�1E3�2��դ�V\',vf}=��+�C]���!5��!J��o����^%^��o�.|}7�)%�'�@�h:�}�=��P�~9;��_A��ԋ[x�X"�X�J�����I!9����O[����@H��,����Ѹ�L$11a����,����pd҄G��IBN���"@F*G�,�XWg�{(,��܌6�y�t���Z-	�$�+��_�u]����Q��J�af�n�b�rb����Kj���̯�f��9V�"� ����@?�À֚��Nf$�)��03Z�u���{8���&ie�=D��_��H�S��Ey�6fF���A��/6�#qw�/g������z���p�l�ĺ�:���rPkYC�@asÝ�Ƥd�hξ`�7CK���O����<j�A2��Vd72�x�&o���k˪�%h�U�S���4.�[`#��&�z��T���*¦�H�z��[@c�j<.�pXr�}�b,	��������mB)zV��.�D��{Ǆ(.�C%=8��Wn9y-�����`Z�����eZ���gosh��R�MZ��!ۀ7�Z��;�$⪞J䗳kO�f����]QPJ��C𰴴T���WI��'�$���Cq+�	11øp�>��9�<���J�-ƓP]�VA�ׂ��W�U�}N�Q'�l�h�NXeS.��"��yC�@Y�?ہq\��f?�z������ET1�.o;k1Ђ�>CY5Ը�W�;V�-�O�<F�W�31�ҿh�2����}�����w��V��Ob��^�$��I7�����Dk��ܲn��د�DVn��n���K8W�&���w�Wހ�<⽯55�Ѽn\�R�߭��O+���B(k��k���r�D�-����)B5Y���G�[i���z�O߄3�p1ڡ����E�YMm%�VTQ8b����X�B*�� ;����I����,�Be^�'z�i����l����al�#��<�.흃�b����q����
�r(�t2t�3���Ca%[G�ض}ݍ��
.!yG�u=#�]����~X)��l��.o�U׊�B�3��S�.e�H�Npr��A��$�O�/Oo�K���P���	G���=�����xd2��[��U)A����C�2��e\���À3������$z��X�:q��d�P^b��t� ��G�f���V"�d��#�ә�+ԔP�)o����K���7�k�"�A��~�zACS���$ho�3�q���.~��KjX~/M��km�E�pޣwuؤ��c�W�V\0u��� ��IؿV>��V��SCp�+��2ـ�᰺G���BmGt�V���ŧ�,��&nk/rQۍh?8�J��S8�����ʋ�9m�� ���D�~"�l��E�E,�~R�c�e�H�ץ�Շ,�ʺ<4B�.#��M��&ɻI�3����Z���v�b�b�c$	4e�eR���5��}�m���~6Ĕ���^�i_���O��Ж��fb�&7y����c�g��$z�Ľ�ޏz��`����#�ȐcCLl�5N���ࣻ����bbV1��Lz��ڲ@R��3�1s[��m9�C�k+e?Sǜۈp�OL"�A"vS��2u�ܘ�D:� ���|.$��䤱?�&�B�L��mMNX/6��2F��ߊ����@5ι/���Ǡ�qz�S`9S�C D;FS���z��&fӜi?��|�-��?�
��m.BUg�h��AB�˃=�q�]x�tG��T�����q�\�I���e��c�i�xz�lgP��|���ݫ������� ��D��s�F��>z�7��Czl����`�&N8�','g�6�"�2��wb��;�hX.z��2V�|H��������>�H�A�h��]$����cF!CL�0��G��,Ѝ��^`�Wel�w?�'N�	[f�s�0C�$�rK�� D@�|Z�i7�9��8�ϫH)�%��a����A"f���B�4r��"��Ldm�=��OT�zf�qĬ,c���}�"�ħ��~3�x�
A�,����Z�U9���.��b?��SH�E<�h���"\��8�%���.�i$#p�*�"��
�E�!�sz�ԣ��	�=���d1QO�W��#�uςl�S�=��Y<�.D2���ȰnO{a�t͖���o�-\b�    IEND�B`�PK   �A�XP��/�  ǽ  /   images/f42d805d-3c79-4d19-85d7-77e6ec425ca7.png\�T����"  "%�R"��%�]�J7�ҝRҭtww�tI���<��]wݽ�Y.����;o<����U�GA�C���A��Q���u��y���s}X��y�($����������H����,{;)�z0�VP,~gN��,khm�l*S�6f��}D!3ܤ��VR�q{�Y\ÑV�]'A���fӵ4�ϓ��q�K����y���q�=~<I�����ӗ!hG{��%�M?�ă���w-&O���;z+8��Q���f���~O�&��D���?��e�yJ�@�-B�����z%1�����>&]���b��bp��W�	�H(a�o��d��-���Q�+4�R\�xWe���*.4�����oq�`��F8��c�L{p��ڢ��}
sR��z�S�!�����w�
^~&�*]��R�\H��sݐq�g�A�*�{��p���_���tcd�=㬖T[`��e�b�^Y0>Y��҆�R�L���y��up������$:�+􇇇�q2o��h�ۮ|�6 +ݐ����%T��0+�U����"���7��\��A����'��KF�R���������Jy ��a��υ�;�f��J;��	}|��j�b�i�]�|$1�\��s� i��~b�ͤ=,
�Ȁ��I>��[$�m��-"�c�V��g�~���'�����K��k>:,��.�"C����H��3�_$2^.<�U��)�	W����
ٟ?���*ȥI��+̕b����b�
�Tm&��J�](H��7{���w�xc��%"ҽ�Q�Ύ���<���Ͳ��kNtttfף%���qj�ES���.���8��a���A�Oԧ	�XH�?�����K���s� ȸ4w0��.��\�g�?��涉�Ȃ�E�L��/ڿ�q��1�w�0��ßj0�������@*����8�����E{gm�R���AY%ߣ���<,�QO}�o���04��=����_/��W��"BB�N�l��0�\@0~�h�U&H$�=��?�W��� u���YLAL$��Sh�,�٩�ha4b>�<P%oɁ�@����S����ez�R��M�/6��C�i.f�����oӳ�������S�ae*���r�|%�|%�MV��0"u�T����B�l���2w�$����u?I.�ꟆU�nn80�����00x��0�������CnbȚ	3y�6��7P�_,��
D*��{y��?�%���&PRVN�!��d-O��6�_d�����ѫD��,��V��c�݃�k˩�$^����96�
Ll_Q��z���)�����%��'.�7�ٓ����>�$g�_�1vm����
	B�^��z�t	
��;"$��UU����.���f�B�փ.��'�����뙓 �vHOW��3� ��S/
�����?vW7��KF<jF��Z�G��p�����V��GF�;�uu-7K�Ɉ�(!�a]�"���T�OM��<7�DE�待6���V�!�iJ�%9�f��f�����S�?2ޤ��CNS��m��^�?=�b��vjwZe����R>(���/�%�SF�'�g��a��渶�0n�C6�l���_����o���ͽX"%ُ�
����cka��,x�|t�|rE)Q���;��Ի�I��_[���W1Նp���eK�w5���b��k!0TW;O�/:"��M���{c�;�_�|E$��E���+�eE���K�k6��	+7�-��I�t�S
�^�r#^���Hw�k�����!��#�#�k�K%%�<\����D-���M�=	�F�dq�8�455[|�$��42�˖�p���c�٢Q��X^E��\�:��祺���Ĩ�sh��7n���sj���i(2T�E*aY���;�����LoD�Ă��G�����=S'owk���K-x_����>I�����D���Z���Ͽj9��!CO�7���{�K���dvu�o�W��aA�sbaqS)�1K�"�w�Q�ӳ���,}9*�΀���4[(���8��`��}�慀!.�?�XT==��0�*T6Ư�"�ڃΏ[���l%E�R'fH�p���E�� 4a������ײ�|�b1�c����aID��9wf��X��Ku�0���d�0��,^�c?_*��+l"�.�������k���Թ����ܽG
u.6%��M���
br��O$�N�?�?�bi���ܛ�\~�u1t`�0�AS=���~��3��e>z�����������uR�@�h�|Y�+�9�qM47��B���F8��&��O���\�p�}����uJ�y�H�k82z��_��9�"�5��`-��|&r�LS�Q��+%BŠrV,*����#om�.ל� W,�}9�@�p�H�����'����P�6�"z�6���?����aF#3��|8��?N�~{��;6��K���14��p��% ���8[r��N�Ȧ�B/��W)���e��ckm����"6I��ߺhwFDD�WEB��(qM$2)�X��E�/��$j?0T:9�TU��0�||��M��sC����(e����jZxU׷Q�
�}��i����D�۩a�� p��	�SvG�'<��ƾ�ãV����	MM︤е��Xp>��%G���*ӕo�"]�b���Õ�P��el�{Ԙ�� @2}�HI�X֦����ݱ11~7�;w�����YR���q�����&�����hn��,��Fg�؇V�S�^���>��.���4�榤}��������Ot�"+~j����"�%�`����W�
}m�?eT���u͝�_�Z&L�F��CDL�����9A*pkkˏq�pq�⡮���?�xW�I�v�SR�S:���J R�U��0�-�u�T��!c\�W@;Gj�p�Ic�tdd^��6��H?�v���_c����Q�C�� _��\mh�,,ts=��D=�T��_��+���_+��1��"�.5Vѩ�0�9�HW�
������NŰiL]��㝳��ԓ߆T�b-N4�X�!�ѥ�*7 N8h��׹��:���0�OOˤ�_EtَD�b��ţ|b'�
ޞ���QȐc�7�bq�b2_Ǡ1Nhc�1Kp�,�P�Ģ���o���F��� R��r�eU���mWa���Ƨ"�9��+k��uZ$�*6�Ud��Y�̪�a���W��b���K���t�<iק�)Y2�p����Z{[l���;=R�Kţ;|6��x�Â>��&�h��L]Q��ȒQ��W��\�E�����8>�A�����,`�E�� �y��7����YQ,�˧6&~qk/^���m�(�M�X��O������_�.s�E��L�n��PBv�l#����c��J�&�<������,������>ߧY%t���T�>�K������&t9
��چnA;���	����"����?]p+��hm!]��r�?_I@9u��g
G��\#��Z:O��0����5V?_|H��
v�x�&j�\ϥ�W~��s���z�ֻ�!����	Ve[�Su��梦���{����z��l���kr�V���s:����G�M,�<t����ю�a<`%
�g8�/�lG���'���n��.���y�y�0@�Ȇ|A��[���_cbR��"�pj�;�=iD��YN�Uv�����a|?<��1�+���ĥCA-�c�ig������D�DDV1�-���DMArѿ�_�m*���������²1X�M����X�t_����05��0~Ã��<��m�=;�M|�1y���ъ��݇fB���f�R%�Ye��4�i�S#�I�{�y��{���ȗw�#3U��~�#&���ԉ�ls�S�����Jb!v�Ϋڨd�{|��a��b<���0
��o���ajb������n��
K��gr8_f��/<��W|���V��20�"O5�T!6i[m��Yk|�Jhy���H!x�%�A1|*�v�C���h�h|j޿U>��Z���'��[��v+�bnv��@S����Q.J|<Mn�";�o��Y�|�[�o�h&ȩU��Tc�p,p�Z��ҼS9|�B�e�:=S�e�o^|�Or:;;v��I^��K�5^����.�͐�ު`�p����E>�á	E^�a���0~7�A}�e5�����.��\�dHu�3����ol��b����1tl��I��?��ҿc�ś�BQ�1(����"Y(��W�����=�z���7�Y��mN_5{�z�,
&�������9�\��і���-1$�ez�M�o���E��{�֎Kߞ��b��s$�J4�v�?=ɀ�N�:���Ԋh�J����Ս>N)�CJ�FW�%���iq�t�0/Z����0��X_b�ǂ��4����S��J(DG1ĭz��.-��ѧk�qpK(1Q����q�]X	�"�C��vf���*�Dy�`�����ǳ�!�-ň���C�/oq`��Ia��f�K��4�s�:�^7a:"���\�+{g���j�G�3z��A��+?������h��M(C��v��[�NP-&���{�e��O���q�!�9���>��>4�WX	*I7�;��݆���V�5��� H�*N��zB�I��}�Z��*�n�ӣ^fk��22�;�iqf���O�n�%����$B_&��W�������V>���o�Ҡb�W�&Xߙ6+I�RM(w�(A�`'}7���t+�sC;���x�������.S7R����eQ��f�&('�
�� J�&����FM
< ����U,|Θ�JM�_;�p;�;���N_�^T֩K�b�{AU��6�1�.5W|�����|��WX?��՗�|�N��y�lyk�V�����w���H�&��W����VS6C�+_F�}���5�ɪ>m'�Uźi��9X:(rJ)�����w?��Qu��!>T6�.�DsTr.jvt�|���k�C����\���r��~v����.�B�� �G�i�xJG��˗<3�vv�F�A�B賜a"Ga�_��ε4c��ɽ�:6�W�M�˵��B9�q������~=M�n��8�a���������[�P��
���uh�����A���g��vF��zk�/[��aM�������L�sR�ӏ�Rԯf�T0wE�3�Ԣ'�jl�;�0ˊ�=�6�3AuH��������0�7��F���XKX|E9#).'��FK��
װ}S���nǂ��,��jo`�Q��l+*�f�N��ox��x<U�����Y'��2�P��sɄ*��]SַHf�t_�!ى"B+ђ� t*� ����W������7p�_K�UU��Ⱦ;
�<MWZ�1�r�'���$��R�E����1D�C=�Yi1����U���_nC���	�d޲��?�h���:6�QJ8�vB`Y�CjP'8�̋���%�D<��2	������:V�`��<�#�<��P<uK!�$�Ԍ-��ѫ��@>@�v:��Z��n���a�̆ONl�_|��Ϭe�2��BX2Spn	z8H�P:��r��N@C/V;�R��9-S���|�W����*	�m���
��9���!�^<E��#9�%�!�qn�Ÿ6&�4zU]7K�yQ0��ͱ��?n}^�WW3O,�K���7&"�S�#�>�«���p6�LN���/�2Ďywtq���$x���S�������zh���@�ʾ��Ef�S�Wt��z�e�A䳴h��F��*���a�)(��
�
�mT&��M�o왧8������n�Aɍ8{M�6�Y[�u�Oq�ᵃ�A�׌�ڴ��RMK�-I��m���ϘõdT[��SW����t���*N�-�ҋϲ;��%	ג741[�y��h�"N�,�_P󣄗�V`:��hS�xQ����j�k9��3bCHԓ�{Oi��#{��dm�O��	N�<�m59զb��#"����ܵ�q�[g�x>�M66��ZC�h6��?]�K�X��c��ta�p4{Le1e�i3�<�~�8{���g�,
"H��Z-[��+*�3\��1���~/�s��K��Z�#qܢ��&�����~����,tO��
�0cبu/�(�U9��Y����Z8���һGBԭ�g�v`��$M 	/Ơ�2�K������N�ևr�ބ�1�ī�,�k6��g�^������c��%x�//EX�{!h��t����;
01��,P�<����.p/|� g�t��q�)���od��em_Y�'�3l?�熍���4�pm&cĘ!N��3G�ێ�����s�j�3�47���~�B`Ts�b,ω��-����s|l-��r���X�غ7:�G!#��n.y�8���)wSj��C�_�*{�1Jʟ��Nn83�sԼzы�ɕ��F��Z^���K��Q}�i�[  �l�$/m��D)�HH�YZ8�}��]~3�=�"
=@�q�����L2e��PF&�cr9q<ҋ��d���-T���O�����)Y��0a�g�ܟs}ρj��`�!&�mX~��u}s�"�M��n��#ꀺ*���}y������s��I�>%J���d�_#�=�a%oV5������>�P(�ph�˙?��K�rVm�/�Q�g�2?�e��gɏ
���xk��f�N~]�����hE��2*:XF))9#��p���bz�3�|�~Z����16���`uLL�_�����}��H��^���L�}��/�!Oo�?�Z���n�����kG�_qW�}�V|��y^]���t��Q֍A ��領>{I�P�c�&�"r��,�R�S�{�=^��?^��q��[fy?���k\���r�|��F�]�ߘ֤S�_z�6�h��5���S�v�qYzM��o�5��}k�noǙ���Y<�C�ƕ����/;�r�T���Զ������\9�9����}nH9^y�O{=à�'e G��|s�iɴ����M��f�_�X���a��m����r!.d��C£a�[x�Pռn���[�b<���L{���Oq�U�:��Lz��F�U�9�$�:�m��#��M���Q���޸Oدm��>n���[j��Q����k�f���6cbZ9�}CU�:�s�vpJ ������s���oƄ+=y���W�%Za��<Z��ڹ�/2Ƒ�K=�^�������gJ�V���A��v�����K�#�ߦP�Pf���p#U��.2�ϛ%n�TsNy�v��~ͯ�w��=�f[�p�<���>S�١s�|	I�&ˡ�P�	�[�\u$5��1߫�;5�������}��;�l� ���S�jGؙEzI���F��2M��s�7�9�/�d�BBr"bƞD�A�Tn�V� �}��t����s�)�
r���K���F�����H��hDov$ټ�,]l��>�9�+۠����z}�n�H�ȋ
��ʈ-j�"���qAl'��%gA0�ϸ���_���K�tt�_;K�*ѣ0�dh�2X�ęs�n#܉|/7�@ =
��
&��G�t^��:������Pa.&s�:F%!]�m;��pc�[G�'&�\�`���J�B�X[ִ�7ϲ�^�H��+}l��U���;\��rg�w2��[<�b�;jo���=ryCg�-���d;�q����)�|V-8hޥ�C�,�XVXH�zG��I�.k�4��{��Cw��IG�篫qK$�RT���oȴ��%X�u�2�BE�#!R���k�J\{@��p�	����(��j�9�|���G����Ifz���V�곾��ϒ:�Z5��n���V�܏]�ֵ�_�a�����lN�f+�d)�����(�o����C�;��Ȭ�0���k�	��_:&�lcH��ly��:�~Cn0�޶H
���\L ǁ���b( vlG-�w��,�������_�<�����m2�;���}�#C�v?���9�K;6od�mH"ÅV_	[��A�|��l��'iD|&mn>S��j޺�����A@��M-ox��v2��߭0���v	���� Z�՜7�dnP�7�|r\
e���f�F���I�>�Ev"Z�$�e��9�O�8^[c@0��0�UU�l򎸟�"����������酕ge�/�Xj�q�N����X=;#�����rP9s��=
��~F�U���q�dd��Ё��o�����v����ԠayRjU�[X,Q�D@�O�Bd�=��l�fF��u#�� 6O)��%���_c+4�-�E>qڋm�������8� <Hd�߼ϕ�Q."q� P�s�pG�	�#̇�wq�x,�Oi0Ϻ��7Bf|ۺ����*Z��+�eQU�";[�=���f;�3���-< �E���p����( Ԋ�E��J�]����ec]�B&�++6D�d@n�p�ĄH�V/����9`m��˕�F������hkk�벽@���<�
ݢ���aT�0.a~���V�"����E��iPnp	�ǭ��beU��+���ddH/��I���?K��N⯢I����DU�eR,*���8(�H�j�

&���~�c���՜��7s-^,3[��6[s7�h�,h�5J�9��
���k�*N�����3�P��)��C��`�nYD������w�CZG��jk3�j�������{Wb�4��`I����B�Vz��i�����5����G�D�t1J���$�f�5w���M|v08:|�����t�7��p�A�R'�h�d�B���(AG	����-��-\�FA�b��j@BԵ	
4�˝�V"x`kB��]��>)��;A���0��A߶DZ��t�@C@i�C�_�*��mmS離��i*��-���qI��NS��Qx�����>�TIB4EC%q
��=r]>&j��Oh<�u)c3V�lb5�S4#:~Q���}�F%���R��u�DQfG�Ǻ�B�<�c��	�1��^|�r�v�X��w�3*��V�����BPN��<fY��=d���U���S�1��t�K��� �Q�l��J����h-%�CWH�~!�*n��v̞��ݶ���MP�ٓ���h�i��]�����Mg�ITÈ1#XX|v���j��lE�r���,L�Y����6���v�g�������D��bK���J\�M3���q�H�~a��Rx߾$�3Z��Pm�slӂ�O x��G#����u���A�L�����F �C 0�*����� �]�.ߋ���E�E�:]e���R���y{�2��Όߓ��x._�z�At�f�|������'��!��/�%4<����-S��A%��冽y�R@�d�rL��5��E��BlR`	�|��5R�^�7��l�1�w)Ӡb}�0���GD�}ng �Ɣnӧi�F�l��H<��j�R d��$R0�?)t�1�=O���7^�╍�2k"��џ<�L�ݿ�Mk.o\�Y[.��jY*������a�M�M2ׅ�$�~!�	���0�Gy����]�br%/�|��^;��(�� &^�<��1��p����Z4�`��F6�T7�k��G#��p"�D QFz��j[�z7�G��n�cpS\� ����&^� ���aM��k�D��v*V�@�mù�("	k���BS���od���q_?��9획����OP�B�I��+rY�(�l�:�����zL�"O3�*����qZ|��u�/f=��`�b��@æ� #q�]k�?a�)~�򶱄�h0j՝gǮ�#vIdShIs,���˗����A�PDz$�~�%�����p�-�C��G�����w~Hbn"+G"$�w���_k ��[d˻�����a`l�����_!�����Gf~0�/g��[���	AT(�jú�(�U�l��g4��ul���+��^y]֑ex5��nLpǐ \"�.���u�RYLA�, T�3.݆��Z�q5(F>(���:�|@��ٵ��}��[���LN���
�g���	hh�ҳ��t(�T�HI�)9Wq�����ק��IP����V��ܡ!!���!:,�1�	�B�zj6�^ ��c���I4��x��$�4���O�k��JG���@ރ���>�K���ӈʅ��B;u��{
/����S2���B/���{��	_n���}�����
�d�T��ٳ��?4�@a���]��*�(������O���T�ȑ��`�HU\=yr��Z�X��an��CdD΂�����4��5�#J�5C����D�48I�]r�n��r�x,�
u �4�w4x��"�X��S��*m4W8- ��$��+����}^�.}���"��l��S�M��pP�N���H��+�B�VbKq��������Ҕ������n�.��R�b��V2@G��=~�a �\-�BA���b0��>��� 1���5����A�����sC1��� �D�;�7_ r?m�4��~����7H}fx
���~��Z���~M��9��.�*�nk�x �5;�&�y��*����+�`�T����K.��oD��x�7$�ut`==á�b��R����t6P��Ǐ�B����q��]��'_k�R^����1Mz��z��Qf)��E"����4��C0C�>�<��yE!���rK`Y*�=�$^����T6�Xɗ;�%�JA[Ԩ�[mH�m��Ph"�-�$ݗ<�pt�)H=)=:�d𨎿N
1��߯ 0�Ej��\�팷q�q����s��p��.�~�b�y`Aa[4�J������"Te�CP�����"�9~���=��g��9Y��B��[&��Π����e�o�����-�3���ǳǾ�h�UE���9�
�ʐis�Z)�#�-h�W�� '��]2D���&���Gƪ %�02sr$��(i�d\�
�1ެ5����(���X���ڟ$���T�li���X
�R ��"�o�l�FrPQ��m>\�MW����l�cn��e6YT����_I��8�����ⴊ�:���)t�tj��"2�J�ۗ�ǃ���������Hl�K+~@΃�Wh}�Wa�<�4 ۿ�ݲ�3i�"�C'*�DT�^i.ܱvۯ���>�0�B ���z����=��:C嗣&�&>��C$iy��>�<#;x�vwե����@�]x��#���<孷���j�x������f� zX�S�aB�&u �z�!�V*�$ UO��b�X�Vf/�l���%�alBF����騜U��gi���>4�kjj��Q~92�ߒ���HT2�e�.�X����# J�s��y�l@�4�. ��4k�&��>hd:� ��6H��e����h&��c�T��b�9��t;#{���#��y^J$n�h���z����J�uȍ_ݠL[k5�e��qH&zn/����A�|�����������<��a>�ջ�l�f�}��py�.l���R���j����_8XW>!?��$��i����s�)Զ�u�+o����6 N	�s���ɀNl����l�jP�K3��Zt�TPnj��g��9G덊@e�(x��[2-�HY�9�Q:�I瘠��:1ǫ]�G��0T1�T�z+��zf�鿻�4��٫8��K�~`�F
F/�0!"g��D�����}�5��Kr���3X��	�2��uv�趆��S9��A��Q��Ȅb�L'l�d���~�]Ҽ�t3�~��O���.�>H���>9�Z�j���l���c��l���؛zq3�O����f��o�cي(+�~��gVB��2�K�)\d~�HHA���|�T�%^
0g`G�Ĵ�C,��B����[d��e��w����w��7���1mh�2��f(���Y��m��xs$����9�lr2��-��!f�!7 l��I����N
D�ٽl�7�K�Φ������oV��� �<�.�*@0�{��i�E�����\K�meߗJ����]��.	������?RPHHIHII�ʯu=D�XMՇ��ݑ���A;a��!�ZG����%Wi*�;/l_֐R԰7 *$OE1O�A� 3�&@M�
{�G4sds�]�a�VE���
������l��� �>�Oh��eyPJ]��]��Q[]�,��o��b��v��<:e�-W�Fɚ]��[�a�Ҹ9[� ֪�=��Oz4#�l�lRX0�K�1� ��z,�4ğr� h�V��� ۏ�"�-��v7)�Y��zRH>`+~�wfO��A��#*_|�7��wbc�I%�"�h^`5Qv�{�б�����8�e}����׸#h�/:����t냆�ҲI(p���k'�&�^-���H��<��}o'��S�t˟tuu-I�ɽ�ɋ�P��@��v<C�b���8�j��d���ː���w�j�4��ٿ�L�I���m0$;W/�1�@
A�V�p>2<,��H+<-�Gl��hM�'�f�)��b��N���#4m���8����B|���K&��t�8�"� 9�L}� =�i����+�b4���\*߫�]̙;������h�ɐic� f���\H���0~#���:��[Da�9�hSq(�Ua1��R����1����M}��@�5g�&� ��m���'<���rn���oR�#��6RZ�룠9�!Sex�p�C�[hwh��UX85'&���'?�����$���:x��vҐ݆�mG��o�H�|E���"��X��~��l�``�@S�����h�X��΀K�$Z��s�X@���U�H��br�����E0/!H �`h�3���a�ێ��O�j(�P��%6O��IE����J�� �0�p�n��u&�Ā���*�}
H��_ł+!�m��݀��*�c�@�+�7�����l��X6˭<�;M��$�n;�e�x�Z��g���ԧ��Il�+�F�m]rh�� 4C@AF����a��6~8
�#`f@�7�)\0���4���<�P �$��X狈^��a��� ;��n�"�l���-�yy��G�dn��� �-)�~�r�x� ^��?ˬ�a�i ��Ѐ���L�138����4�����j�Ρy�l�h^��������	�J��6��Hb��!���`F��i����W�7E(��Rm>��� ���^d9�p(wt䙙~�LGճ�d���	A��ܮ�꽏�����{�;mp�6l�R�1���2��_{e�Jv���(���{ ,�U���!����)�X!��ܚ�(;�~�2!
�����Iyq�E��ݍX�A���C�sw��\T�d����~���9����5�)�l`��90����כMX��[���r����"�#ض̆��r{:����^��z8��Z]�r>��|�
���J��z���ɝ�H���������_�X�x�p���>V�3q�S�WP�T��S�����v����L��f���wu.��V�{�v� a��������g�L���gVi{��,�X����9]K1v�����κ��l,���:��.ju��d��&�Ϟ,2���]!���i�.R�U�i�B;�mFf`�+񽮸ѝ�u��q���Fh�c1N�n�Ϲ|;?���b�i�n}�	���,c����<��O�$��|�5�ި:86. K��I\Q6�yc	��o�r�(hIƅ��A���W�����}}�㥠=.���������m�M�
?���;?^��U�G�~QR�����Ix��	�[���+�_c���8!p�9����y_����cp�j}��p�PU��if������4}�������y\-X~���Q���@�ɝ���+���_j-���#�.R�о�[mkݶ���P����G߉cU�dBǎ�����t~*�_ʨ����o9��M�� �g��r�w���5S�xd�M�����C�zǫ�A��k[��w�H�Fļ�h�Iv2�^�U�+�Ľ����^��00���k�׉)z�F�UI��F�=Ӷ�׍hw�=���\��5dw�v����Q,���r�����;)���� ���2���i[�E{�|;�5^�����9�)�U�-��}&ZS��k�z��樿U^�~�dp�d�r4��u{CJĞ���v��nG����K�����:���@�s�{G7�:���v����ކTW[+�����Qu�[t�I�jG�s>�X�ٮ��8�hEn�~�pGl}Y�_�T<�{�~��\{Y�N�&{�� ����dx���Hq|��w�_�mџW�OZ��%�=y/%�;����W]t:���ӕR�ΰL|�'��P���r#�-F����5u��7Ew{A����˖�� ��yΆ蔲�k�b��}�xû�����Ҏ)��\s�q������ֻ�ޮ}7������:��'Qt�V�7�9WB�O��W��s�.��Km4j����lfD=�MR�6j_��16�-���[�v��7�ٵ&>1U.{��T��AY��u��ߛ�%�h3j+�������'%2��:��X����kk�����KB�2�}s�f���������'k셣k�4q?�8���J�l�%����*4���6��aN���6�P��<wĮ�� *����*7`��$,u~�p�&��=���B��/�;"}򑢵����*=�{�|ԅg#�Ѱ��-���%�$�H<ߓ9!�fd߳.ץ�Y�fd�W�$s{J��AM&	pG>>4W��p��k�DG�l"nsE�8����f�M���3È�' ::����!�zafn!p U.�������f
�=, �+y�e*zW�g zqc4`!O�Gs{��67G����z�&-��r^J���+�$ex݃� 6�_��;�|�}|��wW5p���?�;��+\Q�h��K��L�N�|��滸�5��`!�޾ߴ���d����l�8�V�{����W,�]]��u�����(*	Z�o��NQ�9�/�g��6S�ÌA ;�fM��3$`W��\=XhQ1B��m{�=�:���$z_\i�{k�E-�N�ɣ�����,��:������L����*��E��;׾Q	�� ��(�8(�G<RXI-�S��ߒ�6����4�\��j��|����CL%1�,i��J�sP7	����>�i���R��K����ۻ�M�)�g��p�ܟ$����~�/���z�Fݥ��HV�Cj1@
�]d����V�W�I��l�X�
)�np��\�l�˩��oT�aaV�����	9���Ȣ�~����`9�Ǧ#�M�Ǯ��.BYu����������cH^ �74�g ��eEFwzb��7\R������W �$-��κ�D L���%b��	5���n�&�[Z;)�$1 	��3A".�[?��
s�^;��/�Y�@x�VR�����0;��/CO����1R��
�Sw��8|U?�b��g�O�-!n�p����灒£�?����5��fx��4y�g�Z~��yU��`n���=��x�>��¦�*5M_6�﷿�o�uO8u��OuE5樜>b�94���+�n8c���+R{��|�V~N��j	9~�on��ڃ���ѝ��Jg��(�%����]U��yGc�[9`s^nJ���'	Ԝ��6�t8�Z�ޓN{��6����,*~
�̸�zƛ���P�H.`Dt�vBD��^��DI���S���-O��PVڽ`k���Y��C��Ư#��w��ʮ�u�,�P�jGy��ߏ}��ke�O~�捎�6�5�)�֢����zG���֚�����B�r�"XQ�o��uɅ1fXo��PX]�[��7l��pY��6�I��w�i�z������v��J�%婻oa�E�=]�.�~�G�r�?zJ��4r�H���i�00N���#�,Q#·^n2����6���8 �$B�@�L�}�b�^W��(��}~��dZ���s��Ni"��Od��I����%�8���/O��/糿���?�sK�~w/a�e6��U.�"
���n�ϒ�hh�b�a??�\���h�Q,zG�S��`j���)�~��
Z�y��fѺ+����#ꆸ5�ݤ"������sLWy�������qP'3�T�F䥝����(�4��X�~��l���ğ��t�,�V������]�����W��G�85M�.�F⟠�heU��p��}WUK�?�ե������P�U_[ˌ�v���.b�+n)�n��<�]��?I��$�@�V����uճ�(�?~7��L��uX<�p��7�N3k15Wk�[��Ѿ�k��j}��Z;n�h�?�н��8�e#���+*ԏ���Y��/��N,ե��ȼՈKm�G2KҎ��������3Α��?��SRo x�j&��Y�������1�����\9I������Z����:LPЂ���"�>U���	�*�����O���'�ӛe�y��}�Km���gEX<H�w<n�8c4�eE�H��������M���XZ^�֖���=�3��P�� |��������NI����ZoT�G]��kn�6�t�ܑ�Y�����g7=��^!�늀T��Oq�s�B����$��l��c���/����,R���ѼՓ�]����>��3��(�[a��@܎�/����N	�3�}� -^�h�x~�� �Q	��X�%�/)�D���ao��S����o�y+`p����8��Z�΄]�ُ�؀�:�%���6�.@S7��G��H��.Ȍ���<@�J��e�A�>h�#�'�7�;�ǫ~�<���+Ϭ
_\W�~ݬ����'�~ʓ���l� @dx�uk莑�9=�]�v=sH�����m�ĺ�%�\����4w�Oy����g]xz��48��`�[�nI9��z
,��׮�]{�h��l����o���v�����޿�~�ޘ>�^�Mx��i����W%��ȍ~����p��)���%Ĩda�'rh10-M:6i�� cfA�)%5���>� �y _/ ބ��N�o�1�r�dg�o�|V��5"�ܗ��]�k$y�2Y�Ji>�#��A�.6�H���_�]ND�H�~&����@���@X�����T���c6��fܴ�R����\�)�C�l����z�=��QT�\��V_�x�죵����i�\��.�,�f�ڽ���2��"0����&�Um����T�OdL�S��dmMU�Q19��(�c Y�<����<��p��w;��C������bzV����|6z��Z�0H�AW!E,�8O��Q�F����Qƪ�&,P9��9ƠkA5���rG���W�f�r��y�jp*��~�%��CLP��A����|w�����^��+d�C�~�	?%��d���+e�2�I�����o'VL�U�M��W�?��d�]�{�1K�i��J�~8��sᚳ��s����N����h��{�ㇵ�������{�QA%DDZAJ��K��E��`�!DA��`讁�������{b�O�/��Ď{_�u_�ޏ�E�WD��Rx#v�n~�w�I��)��tR�m�}��xFj�tߴz���,�%.�[�@1>�.4~�-��]�g�uY�d��؁���|BYfB��?�,G��{Kf��d��IG6���(g}����"Sީ�t��eyGz��]]�^�~.[AAM�I)g��@k@zԥD�MQ��L��b���c�D�`_w6�U�f�����9�޹�ܪuW�}���4S�"�L#��J�#!Y���r��;>O:���E�%=��i.k���=m�@�1�ː��:46T�@sQNoma�^�M֔��i=�a,��;h�AY�8��M��@��pM�������C@R�j�>qZ�j�$�i�����<h���1x��L�pM�/���?��K�(�^^��T��r~18��~� ��#�HƵm+��F�: #ؑ��0Q�6�P��)���W)&l�_MT��,�0!`kG��^�������w�����i:��,Y�]���D�(�m���I1f�K���|!��"�e��ȝ�	'�WǵU
�r�ɶCЧ�z����@2d�3���BuV�n�}.����]�1T���8Ʃ&k�>���Ī0I���ًY�l���9���wQ�K˔=��-�x[0�6��#w�����KX���_T�f�S���i��#����_�x���(������O�~e���<������7!S�xSd���B]���B�l;/[A�;oWۨ�t��ݢ�����[ߚ7���9>��24$���G��O=��D"�Yyޛ�2kui��b�׶c��?��Iې��yr&��&uT</ ��"�o����7�}.'�j_W;��H�1ez�E�)fd�E��	�͋�)~@'�ǫ���z�Nļ�!j<��"�@�����۩Ǜ�i<[��_�}�J渗��-+��g�"�Q�vIVWF������C����a����W̢�Z�|�&#�p���X���rb�˚�=Å���e�	��'�Q,L;�[�2�_uE>,����}�=�Lg
6yx$��4�$�5k�A�8�|���]����&�,]�c�u�w>����.�~�ъzM��bi¹[��R���d|×'��(ݽ=��䡯�b�����7N�)~�I�$_<�rW�u��划ĸ8��Tt/w%^��N���A��bs�?}�"�	x`�ř ȍ�W�����&yDh�_��:n�����?����2�`��Rx���-G�S�Ǩ�L@�Ȅ��i���p���S��@��j��Fz���Ț�r�P��;��|�w6ў�r�NxkBN<�Z�NtP���$�jvH>�����~���`<!���ne���ځ����@�����]�:!B�1����!�s�m�Y���r���È���mZ�Z_�p}t�ޛ�f���9��"�Ғ\:�$O��pg�>v����k9/��B���E�k��Ne ��(�`v�E�$wt��f^�]=U�Ć�Q�S��g��F�ٳ�y0��ލ���h��1n�
��N��(E���<��7~$����b���g_O/f�N]q�hH[���M̆�# ���� Ͽ���]��>/���%����EAF_����)e&wa]hI|h��eߛ���gKk�J�mׅ'������ќ�%�PO1��g�@��2�J<m?��F�7��t��I0���kLdr�~U)`s�E� Ѩ�{���jIɉ=edXʓ��.��jq�����Ͽ���xH4�ڨ�1��p�V7FO%\�!�E�̑�1r�3`4/h2��������Um��)�R���ߢM�_�}�S��Ҿ��kbN��[�T�>�-/z����ђ'j��x�Axη_��Ʋ��a�a���^V㔳f$�h`��׍�����q%��jT�L�J[d�t|���*�z6'�db�/(�'���d�d���7�`:q�e�R7޽[�ʲ����Ҧ'��N��#m5"9���0���ߠ�\��KzG���G�Q���F��b��Bun��Rq�J��s1'��3z�(8b2���R�`oX��q��
ὴ�k��Ϳ��?o�a��\�3ct�a��Ez�/�P�(4���5�S�7������]�>�V�T�+�Da*腡��̊=N(��&��8<H���Mdޅk)�n�l|{�������{~�����[���y�X>Y%�����Ԉܯ)�I�\'I<�Cwv♩��BN�����b�ĥ�]A��#Rb�6���[0��n^�
��r���@�)tnӛg?�H�{{��I��/ͺ�`T~�ۖ
\ڮ�-W�|r��,핿c�X�哗~!���nS���ܼ+ho6da^���4�#��n~O����K#���`4%��溧�8�Tm��A7փ*�5yFV
[����Y	i�ya>�ˏ�4]A�������Hp��i0�YE�{��,4�ڗHf����LÈ��;,�� �J}+OQn>�gh��xL��X=���{j�+#��ry�]gՎ�rO���f��BF�|Ԍ4��H�li�e���%�;7�cr*��疝I�W�or&�8A���+Ku$;��7�RO�ao��lr�!	�|�d5�몮]y�ѫ��d�C.���;N�'w��l&�v_��{�K��f�S���/����WI��X�r?!=dM���X�i�.�����I^�.Hg�X�9��rY�+�S��T��g��L�wc��EX�MRV:������lr,�.��M���3N��W��t���T劷�/߾Q`
"�%%��S�u|���{b+���/�dz�6ș����ʓ�
�e�T4�J60ٶ�$0F�#Ll�C�\��^a�,1�'tҖ���Reu��mn��mޟz�M��od�7)�klu�~��_�X��4/�������p�D��u\_z���I�W��DX��HWl��rto�o~e�)�lh�96�$?��F�^@����م8/;�ћ��\�k��r�<�m\f�y���'C�*5;�:��7I)����
qtY^�v�X���<�� 'B�1�V��w�{s�e+�x��+��TK֣�v�e��r,<=�$$$�#�C3W��m����^�����J��UD&}��������Ok񬎑����+�!�dU��Zbo3��������U�Ӡ.�@Tп���?��n�������?Y�n�w�i	��pI�q*uv�*��	�l
M.z�"U,l��c�l�}d���6	Q�#QHv6q��.��Y�daN/]%\�k�F���[��:�$�K�����Fn��Yh�b�F&���.�"޽,q��#DOm7�k)���6��Q+�L�(#��(�Hg\y��VE�H�S��'�?ޫ{Sȁ�I�S�F�n/N
��&�Cf�ɷr�]��a�_,U"�^��Z=��r>�<+z%xr�X�5�0&Ȳ�����p_`��.(��o���
���â?��2D������7�V�/�����_�ܸ)o3k�n0�>���W�8�qB�Ιd� ۆz
��	���[o�T�UK�o,��ׇ�v�������W�,eb���W
9X��%�b�aϞ^�"�(�!/}�c��&��M�7.��|n5�?�F-�E;�b\_�*�蚳�5.���p�=�2ȎR�ݝ������z� zk1-�y?�+�E��a}
EC�M�'�n�+^��3����h��hA��ُ���>6#[UR6�9J��D)�19�<&�kC�� ��ti~m�u
��X>�]:�mۏ*��_$6S�9��?���=�k��N�+~���o���*�53W�ޫ8v��L�P�с@,�����h��jج����
`dq��8:�s;�=D/$的<�*�����JTW�y�V�* �-��1�H��29��M��(@;���� ��4]���7��w;v�,	�9��}��p�*<���p���˛K���89�����u���7��I'_Zjn����ʖ��������$+{h����tBI|Lx�ى�r�W���˔�P��$?!]=���MY�F:泰�2�>� ��Du�M�tb�rr�VnKW��S���,ƕlUفD�GS�;۸�&���������5�5�h[H�^Q���O�fMO�-J-(J�ƽ��P@ (p����ξu�V��~5c��/�ˬ���f����v�*w�ᬩS��=���}���?Y�q	��U֗Wg45�P%�Z����]�p?�����Z�~	���i�y#����(�~�y��K��^ڮ,HB��H�9�|?滹���s~W=�m�$����i��Q�]^5z�c��V�'���r�p�^v�5�z������>��)��|��(o'�wR{�o��8��IИ��I�r���ξG����u��ۼ�4�l�0�+��	��eD��=@���V#8w_��?*��_���7��ųr��0�������>�Ye��WTo��x��1��%�� �(�`�z��/sI�D�o�V`U��3N��쌉�u���5���ŹĄ�?�BJ��~���ؕњ�;2��Ns<�Z�y�i���r�_�)r�~��n2�2�SC6�$җ�b�����t������(�ו��0(y�k����덶Z�H�
��'�K~(!��]��-�h�(�I|<�㓟��H�$���{y��j�����-CȄp���[���Ȃ��"�>����SX�\�����N*Q�ȴ����b���[؞�����]c;��I@O�����0�̭�K���Z��&rٍ|�JXc�L���-�<��t���L��������8Zۤ0�y�~��"�Ef�ۼ�xc��r��<�̬�ץ���q-�(��\nc���d��I͟z�4 �8C��篸tH��/�AP>�ii��0�I�SWEw�������j���(	M|��+���})Mr�\\�\q�}��ȝ���d:�{h�V�.�h�cx�#\��b#����|�+zCB�[+Ȼ�>���W�G�u�LT��)��_A��@�|es�n/�cut�:'|���Ǎɺ8�~@���zP�j��ρ����׼�O�b�R�c�����Y����	�o%<{�|&Mwo�B��|�g.d���(6 �9��i�!h;e��KbM�������"�ک>-?����t���Y-�=QQ�4����iN��7�(b P�s��ݺ�����fe٪��h����H��Q��ǎo5�6��^�&�)�� �e*��.���6��OҨ]���0��#b\� �1���*�?̂�1�oS��ϫ�?RB:�.�k��yR��[�s����=��7ys��rj�L<풐6u����zn�>)�SlQ���_�[:����uq����������_�,���eH�TB���.!|3~�������e�SB<h�`?��*X�7��3xD~;{�<�M��M�0�4����/ �qdޟ�ؕ��W:�'��ZIAϙ���hh�����2�"?n/�!#�������Ȅ���>�ގ =�- X�է#u��_EJ���c^�r��wA�	�$ê�>��J2�.)��L������`����l8].�֪��[���7��W�����k!1��v�u���X�=�{_'�X�뷓-C��N����g��
�U6?!�Z��3x�&)��^'�����xFv :�/E]��_k�\�������S��>�9aF`2�Q&i���_�-�o��mR1KS�5Сٝ�	�|����lO����r��Xu���>j;}�����G���tBE��	�hzP�7�@�i����]I�]K��F��̭9�W7��]��3h����}��mKww����SE���Q�w�/ۉqv�\K�b8��è�52��=� �|������Ƹn�w/���hD���	��x	}w$��MG�vko�Ę2m��7L�t���ӿ�Lս;�t�RK�&Å�t	�I_�ʹ�V�i
��������V��x�x�jR�f!��~��C���̇�q��0'�������a+ϳ��})p/���U@
ܽ���<�
b{ �V��-ZB'Y!�w8�v���A"�p�T� �D�w5�+D��g�[��۽�Phཅ`u�Ut���T�'ٯ���- $�K�7)���8B?HĦTﺎ+�
����7��Ueܭ�?$���p���~��r[�W7+m����`�ω���@��4��;�ܚ��8�1�ʅ"��v��^.�/1YAA:�6��|:���

�~������Ns�S��gϺ#`"%�/�� E��r"�v&^��?~�c�_8��,�J�>%��.�q�����Ϝ��]�� Y�-7��^���Zz.WZzl	��ȱ�\�b��è�uC���s&�6�� ��=|�R������@���
r0�lu��IF�?=fb�R�� � WzH��JV:7�E��q�W�&�Rv"v;��;�3����Y^��<�.��(��@�䂇�F]�J����f�?@w��(N���k��2r�_�� +��,�С.�q~о~���V���fN�6�����NG�'ci����VR-`㸫���te�Wg"upɣ��Ke7�ؽ�q"W�,p����ʽ����b}�k�H� ��C����\�����wo�Qf+4��"�-���K;5��tq���c�J�|�l�Q���Y����t*I-H���zO�l+K��h�UB�c���ճg���\<�r�rS��}�H��n	n�U��~����b.g.��je�B�F2b�?��%�n�\�tV��UZ�@tP�Rr�ټ�!1 !b&r���Aů�>;�ܘO=�'�_<��p1�������ݐ!;ܪ�vn��80h�q�m7�����>��!lW��kUk�<̣�b,/v���`��S[�:G+��P���F'w��c <Z.X�f6�`1!wْ��Td�;��O۠}Wp�EC�~U��ݲ��UE��z��7��/�?M�M��El���C����e�� �� �|8��!f\��ʇ�J��aѷ+?����M� ���1U��EXCsপ�����;�e�Q&)}��m>�w>2�q�����C_�P-�5Ir�]�o�I��[�!���!y�ڵ=_iқÛ��w�Ol�VI\��[���&��C]Z�;��=������^С,�à*A��>`�?
����Ʈֱo��^�+�.D]L��ȔM��C�*@���G+�즶�ǒ_�.�O��{}���u)������Y{��(j�c?���u���c�����S1���^���W�ٞC�ղJ"^�6����[�����J�2��z)}`�j�y`a��4!�ck�6�b�]�x�"+{-A��zNr�"�\`2�}u����Z���t�\��k����i������2\����֏.��	�����r���������|��}�b��8xl}��u�
YNԪ��_B7�(<�-��;�^Oc��^�������O!��<uD�C������8��hB�``�R?�Ҭ(@���q�}MHh}�W�δ/띜o�u�U�+I#�� ��>rR#'��#G?q��<G���Kt�ޖգ��8U�����&��^.�C7����H�PT�*����7m�M��X�a��x{�����w��o�IFHl��t;���qd�]
C>-Rg�.ebe;��D�o+N-/OE�m����m�Ȃg''�3��v,��0Q�U%��6���c(lb)�5�ϬXBF	�.Wk��C�!���*A�j��č|P�]=-���^+:�NK�T�#�]�'���q{�d�L� ���VN �����>=��*pc���Dw�o��	��0o#�X��<j��(�A��B����U$0C9F'���ǝ���u�jO�N/���rYyNɑ-\����Z�d
;��V�6^דv������=!�ǝUȔRW._{��t�C�ֵ�/�z����#������Z���{�.���<M��*|��K|Z�ՊƝzI�B�<k`I`���wU�7Cu#3�%P~��@�XZ8"�M&��f:v���7�Τ�;m�������!�u������]2G�I�g���+���E�+j��t$��{*���=ۮ^����@ł`��Y��,�s�@���}�B�� .���������v�nB��5X��Ωg�9��*Gi�{�9fd�zt0[��x�`���ê������ȫ[�X����-�Rv$�Θ
�����_�H0� Y�r�_���X�D��ݻ�Ϟ���(k��Ctө��.�)V��3q�uEʢ�f��y����K�+>����]���SQaR��KQ�t�ʇˍfe)�T}u�]�r���`l�ٕ�����Ӿ��^��ʗ~���㮝a���c��z�xX�,_n�[���ss������A*]���8�x�m����7V�ը���?].�3GBbJ&'��
�MQo�Hh���8�}-�b�n�O3�ʙ
�4�>�G�̀m��g
�.��H�):=)5�c�$L�����j�tS�f�R!P���#w9U��zNlU�V��&�ʖ�/ŧN49�����E��+��;R���nE9f�����H������:�"�5�1M�x��Ѣ�6N�Pf��ߚ0�V\����p;���"ʀz���m�1����_���Y�MY-��{d�H���x2�v�n�m�4�X��s�������-W��n���9e��|�������.T�k�;�O,�[������o��k��z:�?{�m��YXR���<��K�x]�e��eɛ��s��r�u,:̮��)�'#�E��^��J�aųgTd �`�^ǻ���Z����D�y�`��sz�ۣ���g���`�V�"��Gz��ꍼ��̃
a�!����AV�Do�-�j���RPǱ��}���5ŴiJ8X�5t
E��&��t����]�R J&��eka���.���.e,r��X�2RօҴ� �E1)%�+*{�����:��0F��%r2��-	з9�7`��A���6^���f�-��p�$x���:�*�w>Yb��b��"�4J!��30{���L$GTF7\�e�JE��z}g�A,�O��L�f&Vd��s7���/����c�Ў�Ȇ0R���:�2P�y�����7�Z�&�j����
��������i��S�`_%I
xRC����hb�l����~^~N(!�\�|��ߡ1��×��A�^H�>
Q�?
�5ղ�Y����/ 3|�8�
MQj
�?�wS1Ў6��Nme�G�҅]=+�r�.}�d�CE�bQ��������0���/��S�o�񥚡�1R����?cP\"��79Tc���b)�M�k���ٳ#g`�q5�8D{�(��S���Gps(kDF��]U��C6�9�+�&+�ψ�s�k��c��0G`r�U�=D�ִD�^�n'��-\"��?5��>\��0_��N���U�ږ�ls���E��+�K�~/��Ŗ.��O!Ҟ؎snc��K/�]� ώ쿾L ��p>�Y7]�����#�q�f��O��	Ӓ�hJz�e� fW`��*�� ��,����ʟ�D_
^# ����Q�_�m�/�v]�����X�82�Q��~�f�2W�'��^@����������ޜ{u`�:.��i�z6��L��
�w�,��U��!*'��%,����]�\�{>ԋ|w�}�Bޟ�=���9. �ݝ�-Slo�+�3�^V�9B,x���x����d���5z_-K{��lt�	#J#O�ٗ�����e�~4��v9�,B�:k�IW�6����r��k�voل�*A[B^�b��R��v��e�o.����N�QV�B�,T��LF�+��u7S�QU�BnS��ߏ���nɅ4{۔
�=Tƭ+�~u*')�W���ͻ�?�m׉kb��`���+j�yŬ=���r�[���3,/y�+q����F=���T��J���3#!v��(K�m $��If�8���L�E�([J����[+S�����
��8f��޾|��-���_����a�ź�({:�(q��D��h7?)��ЬtR�9��V/�%vcZ8p���Jf�r�O�D��q���m���3���)��;�_��P�U�`鵰�u��n��l�����7�����zUTR�%�?kB&#�gݷ� $;����xX+W�ʗ�AO��//���Xߕ���p���'A��]M�	���~���q���z+���{#^��h�ī�g�����Ɂ;͗�%�� �"*�.S.kXki���Z�1��*w���-ъ鬌��P7��"�U�,p;����h�<-%
j�].4h�<�Qh��- ��SN�T0��Ȥ2csOӴ��V��_�E�z��6S�SH%�>�&�� ^h�ѻOx���ֹ�|�&O����M�`���Ų�Y���߯�w��C�}�be�w�yz�E��"atP!`L��P���Oυ=���~������c���@���R���o�Y	������r���X#�6w/n���D��pL�v��f�8n��I+�fh���9�㉦�鋯�x3we�/���~��\kR�@�<��$�|���g_�+h�ˢֆ���9�g�?�IXQ�R��������1�%������!*�t��_޴�L��}�(�l��'%X���;sBx#�ޝ�^豬�'3��T��/(\���P�K~T-��Y���y������[�X�
��]��߸إk�g�V%�����S��^1X%��W�}��<��M�"B�p�1�s���i�x�h���O0}�c1��{���b���@��Ǳ���6���E\`0d�\)mqF��#�f�������4�����ZǲИX {j��p�@���ecY*덾\�}��<�T����g���[����9aa�y\J��U���(�v�W/k�,lx0�.?�%��|Ų���gMZq����e���0�$$��2e�8"�;"�,+�-�P
������a}{��C8%nr?Z���� JKN�S}h���p0S�������������{�)B�^����HEр�ۗ*f��u_�V}@��x識	�� E3n(����Y|����nj��!l�Q1/Z�z�4~+�|l���4˓��n�qKe�(� �Vd��;��S_���iM�"���v{��=ܬx�:b�g���by�I.�X�n"_��Y��)��?�`�Ih8ǼN�?�#l��i+]�,�,�~�9=���)���b�w����N�?��K�����M��uO�L+�߇���Q�g�:)�(؏�+�>��/1m#)J�t-����iTe�˜:�eӉ����/��Aƹ5��ùF��}�Ug7Q3�z�+ݿ�}1�8�<O^��C[�w�je9��A�y<Z#I�Wr<pTe��B���i҂�ʵ�"�UӖjyZ9���yZʄ������gh1{��{aO��R<ER�c�۶�~�:�����2`+�}����]��HG�Y���ݩu���}Y}&IO��*+{�޸�UbX��x6D�V�ez��"�-�$U��u�0l���l�̛u8���)r�Zس��"j�E� �a�O-����q>�T9�w�>?��@����LL�q���%2��n?��E�FF�a�͋�[�VE@����O�'w0X��KP�0���I�1ο���G����z�I_aծ�����"��2V���g	<K�#þ���޻�|<�ỏ��}�"FV*|�]WT�V�����t=�d+A�O�i�:���$�rƪ��H�=8��h
�����teV�j��pE��fz\�Խ�n��3/0�w�J"��غW4��~�B�eӊ���f"
�����V��p��Ɛ���H�B�#�P��[��>7�����t��x��m;��ن2�ޖ� u/��KBp�)P��,��B{A��5��醑�~��ݛ�oͤ2~$�˸����W2����-��9�cRGö�����@�Zy�~����������'�Ӧd6_#3��ϗ�^o��	Y��=o[�ެ��q�;b��tQ�_��Ɖ}�+��DP���U��	���^M��PСZ2<�k[)��؅'�Y�G�1m�	�y��q*�_zu�=E�N���o���A_\P�1��3e)���=��N�^�.��r>(){~w����`k���ȮJ�YxJjWR�i.���I�f���f��'��VwYs�:ShT]c�;?W��g������������x���`����O��U"v>��`��wr�S�&r �L(��T��f)�o�}��޻5s��/,X|�Yi�(x3�+�JFfωA��S"�}�;r%�g�?]�Hq�Al�hĤ����tjv�q|�P�{�g7/�Ko�,�<e-t{��{$�y��5�����틳�%�YԎ����=mc�ޢ8�#I&�"��?K5�E}dB7<W��C�*����Z�8[��v�3nV�B,���&�Ϥ^�s���ik��*�H��ў���L���+��|#�e`��k$}�}�Ӭ��ìŶ�$J�?r�}iɅ�*��5���������3���_ƈN�\J�]�f�ef�V�P˭��G��`nE�~%DmQ��P8r����ݿO�����$=Z�o�N�MҢ�Q��s�
��^��V��3�_��~NIs�1*�zj>��jى7�W7!�ui�ݘm(�|2����� B�i�[��s��m=����t:F�߫B��⛤��c��L��T3T�ϫ����R�v)m���?���� Ga��f��H׾��ʭ�)��rk�)J�^o�f��:�F�n�	�H���Ӗ�����ػ�Z6�,la_b�D!��ɑ�5Ы��4o��jHGL�*O�0�����S]������>�~��J��+��"��w�Bg���WS-R�Q�0;gY
�P�O�ܻ�Iyz�ZD�z�aQ�����2k֮(��H�=$������Y��p��@�*���/�ػ�v����"{ƾlj�P0������x0iD� ��e*JW�� ���*eZ������ �v��74�ʟ�Q����N��F��g��p���9�<�ߤ��a�ؙ��Q�!���d������C��CC�$ۼ<cb��V%w��y��yK����u��)�Fuǅ ��O�N�n鿅�r��J$��y�Rՙ/���w$]�	���T�%���Q�߂3�+��s����Sz7]���0ePJ��7ir�0a^�Z�{�!�tE`N�5�+���z�@}�I
����5Ǐ�RW�������V7M�����=�Nh-�dİ�_�(N�Z�E}%|L;�
�h��g
�u�GDV��y@�P�v"�7O��9�~0Q�J���N�h�ӴM�B�8��ۖKU2l�~�n?����\xդ"@h
ކ+D����Xh����[.�=��W�7���r��|#��ja
���6������Y=,��4���;i�?�<�w�\��"Mr�s9�Si,"���v��{�M��Il�\o�S�!�N@z��� �V#���/����qj�d�B7�=n�+���극@7t���������;9	���$���(���M���a%�ۨ��Fs�5}���b��4p@8�5 �����귫І���_b�ث}Pm1���]	�0)︪H��׆��?i�D#�Ǘ�
Q��Y0h<�y��Y�)�SQ^` �����-�Gz��pʺ~�$��6Sw�l���1$ +��zE�eN��b�5��mjA3��f[BL�Kw�F7�*jU ����[ډ0U�-�"0�n�B'�ƣf���=�N	́�Y����D�I1�������:������nN��IZl��N
�?�>��Td)� ��/�*;�"��ͫciA��SlՀ����ی��U�*����*MdM�h�� ����7jh��]S���=�ws��+,�3���/�H�N���&��p��p���ti���
��¿|8���f���@�0���>N�
��O��JC�����8�G#fT~��*�	�C�4?�� m�A;�[�)�_F0n�h�!AT�m^��` �t���r'c��I-��2���?~W�jOi��l+ G���J�ݙ�la�m����p�Aİ��j14{�����,͒`�5�~n"���_��i�����1�,J
��6kp��k�_a|O��S7(�N��h�	��BW�������3�z�L;���q�hq1��)�Т��@ZQ�����Y��0��W��ldG�D�A|��5G�]F6Z�?�f�o��t��2c��>U5��>����_��9�-���%)i+�X�OG�O�Z�P��D'��T"��g�����TxM�b8���٨�*��F�<y�hl�.�-�#�9�J����w���_E|III�}�ity���2��T"rJJe---�����/>8��dvS��"-�(�1�iVI����k54��uQ���)Z�s�5���
�;����l��O�����B�0�.�
�z"�0<�Dl�p������y��F�]�wп�����x�Ȓ�4��d��5��q����P��8���`���0�b\Rol���=?+a���X҅ �u(�F?���8�����_
��bV��j���C�9�]E��{j�8�r�q8���GԴ�������W��;���2f:����;��h��ќ����;UQ��<^�����y���4V��#w�!ײ��2��8�,�����G�T۸;)[���	��ꨈ��ƶG�?*"B�2����֢'�Ջ��v�a����Ш3�Z��|�*��������x���S�V���&Ԋɢ�K�����+��F�bX
1�cc:~P�Ѥ�o_�l�v�&d_����^��^��E��PWJ���+�C��Ȑ�!���1����ii����)��B����Y��ֶ����_d0��B�F�0)֘�J�_�5�9�)�
������`p��7�t.��{{U.\ �p�f����H��U�(��G�����*��D)]Y�sz�B��6��[�w~>��ŋ��W�����yP�1��P����+��i�9�Jî���n�8��{.4E��P�ɷ-��>x\`o��j��~��=�N�� B>&8��"@�J~���_�=�I�2-_nn���V�R��Q�`|�x3�eg{�o�"g`p�3��,O�cU�qS��a&�(��P�D^����^��~�ҫ3�L�0���ٙjM�����R��^�I�|��blwW^���������/�x+�\>�z[̵��!��i;���C��Z�B�$��ح>'ҕ2�Mb�k�c�ga��ԙO���5����+X��D�m��}�h��`�Ì�f�M8[a[娠8/
��)�@���q��&��L(��q��(����maj�/=g��V�����Ԣ�s��^���Ȍ��S����_#"Z��#�AĮ� ������?�~}-+h�ͬ��{Tm��,�8[-$$�z��o����в�c�A��!׸}�5fuC�T���O����m��33<��LN�N�s��=��1�� ��#�������p�Y�߳��1�@u��?�d�N���ER�d�睡��s����E�]ǽ7;��ݼ"�/84�����Ν���Ȁ��L.�ɋ�Q��n14Q�v􉍻���ލ+�i�����FY�y�7������w�{�'��ee�g"Us�֚�����[��B�Y_��K���-�p}��]���JIg]��%<��o̊R;gM���4�^*]��s��i���]����W7�p������h�a��j��=s	Q�шg��ޫ�9T�,��b���8}�[T/��$i|T���VIi	��k|w���Z#�M�&Y*���boo$6J:���;7??2""��˩fܑ?I�a:F!;����ffV�+�L��J`}v���]~���!T��]9�T�	ɢRfFƋ���222&\��Ŵe66>�׫�l�lni�`+G�^��f��i�fuS��cbf��eP�(���������ˡq���9�ȱ�Rq˗�H1��o>�����;+��(�x��"�˃[�𸘘�����TTQ����9�rv�k����=7~1nw��2-�t�f�Д����V9����{e�{ص����h�U�2���bhi�i�X�SpgmQ�m�^AᶒV�%+����ohߡ�@��h���z-�3����O�4%'|�'�{c	�$�!��%��-��.��jVP2]y�o���z���@|Lɻ��X�{ff&q3�*�'�J��X���)�U،"�R�Z����������!��T���d�9r� ���7�����(�H�(UQ���g����v]�qq9�B�����eB�-��y���Ř�_r�/�<9�Ⱦf���z�5�����l����/ �ٳ`��@N�q�q���y�{{.y��9 ߽,����Y�V&�_!:�C���x���t%�Ɔ�L�O��fr��ӭQ;�=�noo��`_�{�����$~�+��"(��5�����W�%�����kS�D����۸a�U@E7�����Ł�+;8S{-{t�Q�Q��ji�|)����P4>�i�?��#�z\� ���d���gfeU��K���,��Cxt���~�vj��IQ�kjh�KAЛ���a�gw�b�V��A�
X0��
S�A�sǰz˃ѡcZ��c
�wl*
�E,rd?T�M�Ё()y���1Y�'W��o�f�T��9�����働t^bb�
/�����
����ڕ��^-� R�4����"$��v,@������x���Y�������Ƈ���Kf��K訠?�`�qe2a(����uQ��4-���W��~��������Cu�o�4*6����,���"��J����-<��Ty�p�r�+墬������BL�/W�*�K1
���=�<�?2�#ޫ�l+Y��t���>{D�/6��%ך
��zV�(?�t��#e�!�B�u�L�5h!�3$�l[�{h]� sM�$el#w��m������4Z���Z����T�0} Y�.��qk������ }��	~P�L1�<AI�uwafc����J?8�P!�=tH�Z'��MC���TUY��>�J����\�2Īƨ��D�	h�_�E~H�
z��ݯ_��dq7T�Օg�>�^@B�룅����?P�ػ�� �����K�?��&��0pY��a@u���,����{�/��Z/�B��>L�mֵ��v�]�.����984����V�B4#�m6�i*�ÔO�p���%�����(Z��$%巶���E��v\������%};I������Dj&}^ ෶X'��+W���vě�<��(����S���L��~��{��1�ˮ�e��W<����dA�*��vrDC�
7|~�� �%�ٽg�_��޷wM�?���/]}u\T]-"�tw�4�H
�)CI*�]"JI�P"%  ��"�tww��w��}����7p�9{?�zֳ�>w��z�u�?g�h�mk~���d�H"Gr�T�?S�YPk�uZ���&����X#Z�av�ve���"����Xw��d�^�:�uu�t��k>̄��
�U��%g�����v_
����]p !f��ى����2��_�?���\��|x.�S�(4=]�C���=���>�%<�
�U(��G?:݁)m*7������vz����|��Eod����2�iXe�#��Zq{ϸ*ٽHHmS�J���N-p�����ЌmM��w:�<��xRE<�|N��j�/�%������U`��*��C(mPߑ_�=���nҶ�����Z�_�!ۄ�/}�"�S	D1	���0��-�B�l�}�at��;�5�J���T�2����QfK�w�C�r��?��}p��g�%�:n��o���h>}���ͽ�X2�Ϛ�j--Mz���f���7�~���r��=��I�583	�Δy�Ejzmgn��Ћ,����|<���Ζp܁��Щ������R�|O��n�f��&�N��n΄k�l�aj�'6h��A��4>"�J�%"#���S�A,r�7��/鴺-y\�''�w�oT��~��E���޾ɼ<�_�?W���!*����/O��%C97y��7|���K����k�~L�҅(e�8m��i���M����r��-�[Ai�$6��k�?]W+M��L���8�/�så=��n}����,u����|��W����E����p�W�i��??Q�/�T6#(��h�ْ�R�JG�;-�����5\�e��ؚHJ���}�7�>V8��!)NlDa�9���3C:�ή�>�/�� � r�@���$�&l�G�ՙTooo�p�ZoW�:C�m��i{�HL�k iw��^b�1o�c�Z
�?��x���92��=U���x����c���P�l�V�tdA��ȝ�$��r�{Mjx����6IQ9�WuurR��~��>������}�S
��`t���!�Hp���A���X��6a���d��H�7�Y�
���$b��y+�����j��D���)��+YLo�Y)!��g����D2w����Q�BF[����/V������t���VO�f��#"���}����8A�T��g�U����#.m�郱�>��@���57��j���Wlͭ�.�6��k�j��ք���o�b�P�Dغi��_�����뀋��J�`�
��*4�N��ъ�:`;o.3R��{�6�Fe���lw�Σ=)�H��1q�yW,���
[�X蠺�+����N���xW�b*��y���h��z�pi����ﺝ�AI�ǳͳԴB'����Mn���n��fx�2U��F�d��I_���Zhq�����*:�#Q4���.パ1�ݭѐ�LQ��)ܜJ���]_�5T��@ 4e�ld	�{���@�?�}I�ؘ��G8ˀ��R������_�� ©���f����h�4�ݓm�����rt���>F�)g�^ (A�BSx �Z��1'��?���ĲM�f��<��VDP�����9��G���?�%)k��r�{�g�(�x�ZS�pKĂ��sC���_�X`�C���ۜ_8��P{���mx�Z&�"�{_�O��5TM����\�`�
�8z^�W��x�0�����l+vrr������b<5�It۪������.��;�}��Z��v�o�\�e���Y[�~+��AXDt~|��fBt�8P�D�6ik�8��<�v�K Vq��T�^�9�z�V��|L��{���d�g�'̿�KtYQ�l��J*�a���ޮ� a��8E�^�B��3 @�� �	�����;L���G��c������gi(���MX�������AT�56�F?qX�z���A��<��%`�3B-y�ż�Q������j��:L���擇:��9�~��z�}�h�ZU���eL=U�{���.��Ff�f��gv���9�6��e:���foD\����CB��f|�N���*���=(O�!�~�>e�c��xQgsp�-Qٓ+,��ǳ|(&�OQR�O��G�ύ���r�q���9)))�' �ń������Y�=��'�:�APf�MBm�P:f���dS*>���6��嶯#��{&��l�L��D�啕� %�+���>�m�:��� ����Ὁ�Y���2s��������VM��Bv�;��Х��"%eeK�7��BAGB�5�	�f..�����L�Ԓ�Nu��u�^�4��gW�������������P̜޲!��Tz�}�ob��+��u�,��9�����:�}dF���g0aL�i��%֬X�ٟ�o�<Bղ��
�����I@F�y^fK�H�, )�V��Pqھ��a�V����-q�Q3�W�m��r)��%=�����#7\K +��94-� !�Jfhm��V4K�����4����'<��C:�m
���B4�J��X]��IJ��/U牚;�kc�d �̒r��X���Ub��̍�i�e�����*�'������F7L��&!��+.�p�yi�= ;$uSY�y�G�*=;j�b���$����2�(�́(�ql�)�����z����L@ 1�ݛ���)G_�����`��~2,�~�S��r��������mB�e�fl�|���Y��MW������fNŌ�2����V��sC��Ĝ��~\1bI�y���C��\��)�"Z%b�F��;oWc�g��#���t*�,�͕D:�H����G�yĮD��W�A�`&ϨO�z��#S�#�������\����W�� �lw����us�_�g����H��i23���9�П���!F�V޿�^��Ʈ����{/�Im��{ҹ�Cs��a�Gv��mZl�7�c5��3Ep�ZdogA��m!����ek�#*B��6|V����Nc��;�ĝ:A�+Zs�Y��p�Ą��	�<`��bdddM[e����m�>��94��T�U�z1��������_�G��x>{~Hʥ��WJ}�;`@iy����~���Ӣ�d����w~����o��X���,p�X���z�IAX���p�痣�?|/ҁq���d��������(��TL�[Ș�`i�6��u��ׇ�V���pݸR�4,��&���a�H!n��ͧp;
�>��2�*��׌

�4�Y�fJ֜�C#_v��Ơ��T�� Q!щm���î�m�*�U��J�-Xs+X��W��ٔ�=�T�4d�Gވ�k�P�Dޒ����(�Gv�=$*Q��tnr?��y�L���dɭ��v��]���k��s��x���׌��l��\C�^�	B��!��d`KPP�N� tXNe�[��M��������}�S�>�|1R�dlt4��w�ߗ�I�ϩp~*{o���Q:�<}|ȳn ��g!c�U}3ө¦&����P;f�ϳ�Hv��6�����A�`�2�3s����^FO�l��}E �6L�~傇������K�~�Sz���1M9$���8� y4��k��Bww���o���ȉ���?�U �[��t��G���e]�2#p�x����S�m<!�	��� �4��'tE�����kmV��;��Q�u`ya3ܝǵY����^�ٱg�lOT��/h/|�<�%��%x1�EQ��N�"a���YU�k͟lt���<��y�`+�c�ː��T�k�����|���USe������	]z�$>4�hfI���"	�W;�"�_����	��Q�j�cD5��������CQ����:b[�r6��r��M�1pw�!���l�a�����[����<�i�� ?V���������[(b8��f]�^�w-���&���Z����3|u��]�WT�����ʈf"%�W9�.t�\i��Ũ��y����oN֗��n�~X_���|ck�������h	�KZ�ռ�n��166P���r�+e9HZ�������:���ubf��?}�MO��3�z#��ж�	%����������
Њ�����e��?��5�O���6��|����#��Xr��EMC���W�7P��5���{"BCS����?)qʮ�$����Z\��@M�@-�����{vE3��gf�gϚ��/��pj*m��\o��K��e�D��i�'�����v��_(;�Ó�׏� ���-T��wQ������>  ]��8���2��nK���Z#Q }�(r��%��rJ��)��|�V�}��	��ѥ��ez;�mS����ώ��w{_�)�7n"����2���j5�sIh��ɯ�|�P�ܕvv�+Y��	���^�����a��Ә�ز<���g�x��SP���́�w4���c��sIa�ج�� -~��*�c�G�Â�Bo����{\&l�ؖ�੝�������V�����]͈�����'n��D��	�ͱ_�""��`���D,�1yr���*>Ni��l�Bڎ�D!�T��05��5�k5/,�Q,����6��D�S@����Q�K\n�p7wq�?dkFpD��ar��4Bd.�P	u������HL��<�T_߀�y&�͑4.�˟�-���ߙ<7ܖL`�滢���Ox��J?xV�HH ;п)è`��{���w��4�+Ft�4(D]����V�wVj��*  ����Ն�'��a-��yԛ�[�#a;;;��� mW	/'��:�� �Ŝk�j(�����d1=:�d�ܷ�[�03$�f�j&��C���3���8^�ޞ�8��ެ���`v\�UM���卽ۓ���pD�~l��g�su瀞4P_W��::fJ(-'�E�F�A�]�/�)����=�������ӝ)<�77�5���iH"u�?�4/8�SΝcd^��� ��uA�q�|s<պ�-��j]dx��ٳ��Uk|���5��d��mҰ�����>0�
�P(l���eb��٬�2���`>a�Ƃ�6qp��R�|T�VHt9���?\gMg���g@�kS�}��|p�G*N.uX�I�H�����Bwq���Kt�a��s^*��*�2
q�Iq)��j���N�$�켼�u�����j��ݽ���=�e����?�~�\b����iļ_%Y���{�y����=A�@dd�s������޴cM�c�h/��H}}}�ggc�������]�����r}����?ha�ꝡq���] ^��a��ެ������5P�ΰC�`�'�@U	t��X�7D��D�Z���~��.fNT"<ѓ�!�@�s���UW}��[9g)�uǺ�r22�����C��C=�zEv��ʽѥN�f���2j��L�� ��o}��g&wu��ֲ�Jo�d�=<�<	e�|)v��ZD�yD{�9"m�
#+��\�r�ϸ�w�
Et����1S6ZT���ڣ����͓�4��DG�R�z*�	D�m�=S�p�%�L3�~��Z�9���)n�< �*�[�T�)�[!����l�ht�>�H����rd�y�&���>A�ޒ�X$@�@%w�zAK�%�h�a���������s4�ڜnh}y	i���/����G��^�]��X��/����2�KV}��8-���Y�RlkYsӪ;2��<����L���Mq�ڿ?������|��t=yX�ˣ�L�7��]&۬�5�Y��5Ȗ����ܸc�ͤ�.����2%$�P�Vi�)f!m�ޚ��~M3�{�1-��ά5�#�]r^#��������D��`�J�X�y�N���A���آVc���qR��8
��c:�Z�P��i������H�9P���>�w�U�Z��_~�}�ts��\DWRj��n�����^2�2���*����4g;��GUp�zw�ߙ1m��}=��ĸx \z=Ǣ������c{ȟާJ�׆���E�*��@C�	����$P/��Bk٤��nkL�4�x��z��q��_������GP< DJ���i#n�i�
����k9���襳?�6�y �"��ōԦ����YN�h%��#�������0�^�_BS�\k�m�6im�("CaҠaa+�,"��	�2�T�,�BS�0�kg�c�
W\$蓙0-��?���;Wnޛ�9}�i��3�'r��uQw����"�\��d4���(�t�D�X݀� ���$9Z,@��&a�0��Hqcr�wE��1@����\�����%j�%b�S���`��%S$-�
���nc��F�}�ހ�ڢ�7h�H'���TY 0�I��N��0ǩ�yq���Ah^��R�5��*�^�:W�IN4,T���!1��}��Lz������E
��
C�R�L��@a������3�³��Z���b[�sO �(i����Bomd���C����9�9e��C��8�k!�W�]̶���K����H����)���ې��BxcU��l���Z\E����
���Mx
s��<b�(�'Q���:�O�c�S�_vH�3;�Q�jA.م�czc>�ﺳx�G�S��V�eAM;eSkQճ���N�"�0U��6ʬ����t�RGE���n�@���8���d�k�eZ"3�����ŝ�{Pf�z#7*��T]�Rf5���
�N�Yd�TzuX��
V�y8�F�.��w�dК��{dkHttt�����j���݀�b�'XX�s1�d�����0��54�It���TהԪ�	��f���g���S�R�ܣ�,�i��+i\����I���ճt�EPÅ?u'���*���ʖ����u�v��ߺL�i�Ԅ�O��ќr��gN�ecv�*�
n$���xR�Y�dr�>�_�"���d�\WMT�J,���i��|��K�·h�Y�c�w��z�	-�z��wM����ch� �k=�g��~"/V$�=��/N;P�E��|�R��tG,�N�@U�X��u{#_��E%�5:sQ���6+].��cU�
vA� �a7>fm���n��~�B����]ה.�!�y��w��w"fMC@��Z|��M�1��޲)�T�����H�1���Oi�g����r*�6��'�O�M�Jw]&�~,��˿h�zΥ�mE�Cz"�B$��������Mn�"��?Mi�â=c�J�fҬ_�n*�p���� `|�jNX��Gv{�摙$q-w����h�[����f��2\L�q�]!%��r1�:�U%� 밧����ˤ(͜P�������w
��s�dz��zf���O�����4VKq3�b-V�N��hߣ,�B�UH,��6i�>`��ט�sL�z!V�RgW���m,M,c
U2|-E�����	�1U�$!U�sŗ�tr�KwK�+�6�Ϸ���ې�cdF'�G��O[$MwiOȫ̬ʴLC�ph���t{"W�""BAy?��^����E/샳%�B�6��=<�	N�=O-�CtJcȉI�+P�n{�{�V��^SI��.��֍3��m�U+"���,5�	N�98o;ɯ,������#��U]��k�h:�2�Vr���^�uO����*�T�R��ˏ_��M� ����\Dzo��E�U�p7jѢ�D�Y�B�g����^��D�J��fO�u����]{"�a�ܴB�~H���MH��jI��뤣آN��4Us�b�f��`��9?4������W��m��4ʇz"�2�����bi�
U5t�9>_��*�b�&h�W��nzR.�:�4D���?F�!�ԛ�V��yo��ĵ/1��$}B����<o�}|�m��:�
�t�Ħ�mJ���b*��O�|��Ut,n�#�?Y���	�L�ɯG&�9�YM~��6�cv�@�B�����z���� ��f�c{��m��Ͷ��170�j�}�OD��O��o\�MplmS�.�勬�o���P6��'{yox�{������(��Z�.�u�z�s?Qd��TW[�N�������p�Bp�q�W��Tv�H/�m�����D22�9ѵ����&Q�X�mBoFs�X��*J ��^I�23ۀ���P��8�z%&��@�\�o���]�_� x�&��G���i�����J6*�w!���1���ә>R�޼mbK��:m�]>�Ҍ^4��:_#	��tC.�����P�db%�*��5���ǥ�`%��B�7�����c�ۯ�̭_?Q�]ŗR� ]���xP����B�߫z"�ˬ"mL����~T�MwII\����9�n^���?F��� ��ݙ�o1�VN�V�6>�B��m��������&�3'5��k�i�왕���4)vmH�
3)���Z�5�g�F�2���+)�+�Ӊ|�3�o8e�Z-�3p���s6J�#&�z�ٖ�B>f�֏�u��gI>fI�SS� ��u&�(�N���s��M��|{�	��HW��_����a�<��0�>w)F)�g��B5�xw|�&�������M�rV:�~O�iv̜�N�;��I	�(E��bTp��p_=��z�iJ���]lؑ��޳�V7�k�����{��#��� '�mJ���F��`�`1؃ׇ7ח���R:��;v�Z�Ab4k�=��6�3�w�~"�L���/�y�f67���ÂB�+&9���{S9�B��{]+3bq��1B�xC�ߏ�cx�˺�ٺ���X
t�
�ܺ��uJJ��L���QyQ�mr.W�*\9��}2��(2�n�w��ݙ
��vcG�_7ڑʿ���D��̢X�U�+I�����_��S�|9�Nd�3J���
~����Z����� a*�$����[(�����$],�~:ř��~|rِ@��O�%Il%�����C�EJ&��B���NBx�)�VS]�DKi~��c(m~�� �Ĉ�9q+'b�$'��ن�-`�	�����d����yS�ǚ�S@�ʽ��c=}S,PB(�5&�^]��1v�_u&���dd�I�i���Ӻ·$!�d�.�q�.�j.���,ۨ�d�U��C�Q��?�q3�Zo`r�0��/�����|��)M��t\��B�c$�.Q.ͦ�d�6i�z|r��<��-څ�-j�~�fe�VUxs�S{B]c�����������\�G��#�1���3�����H#���7F+�=�Lʲ�jl��/�572��\�.7�N������!�ZD[[�?Jw%�'_�!��)0)���>Sb�䎒bJ�����)O&�I�
��c�WrG���,�i^Jh1C�I(�bQ7!�|�F��Z�*h��5��n�����}���w
6K�����s��i�@�'�߽�_�\����'�DQ��D�K�I�JD�xI�<�~4�F��=�7O֑��l{�B�PO;;vdD�,���5�%(v�HapL�M�8�Z��\�}������!����xy<M�R������a�������"*
	X�оNLN~B{��x%��Ww��7pt��(���8
��(`���	��y!7����{�O�~��ǋD��K���멽���$Sin���]��Ck͇�cJ�6� L���rA��c,т}Q�9;�����2�\��t�+���?1��e7/'�����fTr�1����tJ����iE���8�{f���v�]1���c�5��9�)��"\��GıL�'�m������]�M��d�w���{�nO�I�p���d>�������:r�f��1���քK�Nn�ԉ�)�UCib�����,�/��1�Bsw\뉬��%�$AX�V!���cʗa��| �Q�ѯ�!��/)���W|�����L��� ]��w�uO��yWz#�Ƚ����v��VF̊�N��� Z����G�y�X ����g�lX�&O�HR�:p:�ݻ@���O�R�e>rj��)��?���G������*��"��h7�>���R􊨷��/�~��d�UЯ��D��B�Vx�@�G�ٝ��
�@.��]���Lv�Dl��{,,�%������G�!�B�~+I�`���S�wg���uvٸ*������ڃ��9m�he�wL����O'�N��HT�A��8��죞�{�!t�������!k4n9?���,���Z3�À�_�}Ԝ��U��o�?�H�!��$���x��-m��A?�"�ݟ�+ʪɔJ���PK   �A�X�Ӕ  �.     jsons/user_defined.json�Y]o۸�+�_����7�n�)ڤH� AART#ԑ\�n7(���H��4�l�	�}pG�����c������p9է4dy��h�-T�,�NpB��|��G�ã����qbo��*]�E9�89��]��eu��*}Y,�r:��j����ev:�a���Np̐#űGS��cpE	�9���$�}���I�_��{�;�4�X��yeO�AZ�
)d�
oU2+>ø쫫��;�o�Ѳ(��,/����˛I>�M���r:��j��_?+�7��j�j��E�u	3*���E�C9X���r���O�
a��o��q��
����fj]���8�85�uÒ6,�]/�������^XچQ�ga���+�`Y�.{QyUE��~L���Q�oN�_�l��'��(�Q��p�T�Ai��b�6fc���oӊ�������IE���A۔�q�?���mBѸ��~�6���#�w���|׏��(	;��vp�����m��M+B�p�����EX�li�6����'�-�OZ�!Z2����"aM?j�f�HTݏ��X�kǠ�~�6�(�D���m�5b�ڿ���b���"�.��O/�!]"��]�C�d$j?�X�x�HT��Ucc?�������F��_l/��Q���3�!Ǵ��2j�O��{V��P-�utX��j��W�fVԱ�N�M��YbY7|����_��O�����n�u���繛��kU��l���zy�*�b�Y�XVL�^�g(k�aHY�bq��SV��~�J�I��2���O���м�_��;j��`�rpS.�j�V��f�c��r1[.��+�o�RH(k��&E\fi�I���MWV;�N�3HW"�ȥ#�y�Z�3�m^�}�d3�F��:&pdi�!�����R��-ɋ�Ā ˮ���޾�$\LF���cCv��Ӌ�[�h?<2X5��6
�9n�3���#�`	(7;�	�<m��$DPNc�Y���)�,����5�d�ʈ7,!�K�{��E��h�W�'X��5��/^mEםm��T�J��j q�^��������N�
I�.��Y�t��g�L�MQ�뗢w�*��+����_����0�kj0�vԀ��'�Z*!�+�lY�K���,R�9]UPx�
[bN���]�G�-��������_�9��1E��cpE�O����ҕ���)�	����U����|�׃����;���_��qj�j�o�I�3ˌƈ`�!�a�$	ac}�i�E��Q6I*Y�i�3��ma��Q�4V"���M"*%T�ik��d|�N0g�S�G�$��w�$
duoO�DM����+��&}8=��%1��Y?�#���z�cR��ın��q�.�10��
��N����GL���}�����YǥF���ٔB�����5G(�s�����b����3��b@�:Sj��D��sm�l1LQ��)RK�LY{��V�2��ڲV;b
8Y��h�.W�7�SD�~�=�M�%n�_���i�#��N��S�;��7����'ql�T����Ǝ���f���cP��"T��wRy���������ߑ�Z�f@�yL�PJ�y�p +&p�TR�Y����"�U�"+lj8�J�4B�(�=����M;HE��������� �+/}�:GR�B.�M�;b��Y@��Cȸ��	�t�9�=����]:w;xl�:�k���|�k�����g���-��L��32���@7J3�TE��2�gw�ޝ7���˽�H7������z#��4�`��/���K�!�oQK!Z�W��`�c8�K3�����$���t�g�/D�?�^{�,��,����NeY�S\8(�Ő
�:���[����;0����;0���Þ�aW?�PK
   �A�X�2#�  ��                   cirkitFile.jsonPK
   �A�X��_�  >  /               images/17d126d1-8a97-48c5-9cdb-beb53ba7b71c.pngPK
   �A�X�K��]r  ��  /             �.  images/2ad7430d-0d07-4e15-a76a-a5ad941878d2.pngPK
   o�X���Es ?{ /             ��  images/58ea960f-8973-48e4-ae29-a018cd448a26.pngPK
   �A�X+���  D�  /               images/5cebb09a-e86f-4cb2-800e-22da09d26481.pngPK
   �A�X�l��A Ԥ /             [� images/670050b8-4f2c-4603-900e-28b8075f4ca8.pngPK
   o�X<5P�F HL /             �� images/725e652d-7206-4b68-8c1c-12a8993f9b75.pngPK
   �A�XJ���a
    /             �& images/7b1dbb47-bd0f-4b1a-b2fe-3ae5ceef49a5.pngPK
   �A�X`$} [ /             �1 images/a8bb870d-02b9-45f0-bd60-404fdaa8f6ff.pngPK
   �A�X'�Sz�  m  /             ��
 images/b4b7fff7-3733-43f9-86f3-7eaab1c92eea.pngPK
   �A�X$7h�!  �!  /             ?�
 images/c6364832-c854-438f-b38b-75bf2a0cd33f.pngPK
   �A�X�+�s;  z;  /             ��
 images/f3037bb0-f56a-43e4-a2ff-17056f7c669b.pngPK
   �A�XP��/�  ǽ  /             N images/f42d805d-3c79-4d19-85d7-77e6ec425ca7.pngPK
   �A�X�Ӕ  �.               �� jsons/user_defined.jsonPK      �  i�   